magic
tech sky130A
magscale 1 2
timestamp 1672748041
<< viali >>
rect 29929 37417 29963 37451
rect 38209 37417 38243 37451
rect 1777 37213 1811 37247
rect 10517 37213 10551 37247
rect 20269 37213 20303 37247
rect 38025 37213 38059 37247
rect 1593 37077 1627 37111
rect 10609 37077 10643 37111
rect 20085 37077 20119 37111
rect 32321 36873 32355 36907
rect 32505 36737 32539 36771
rect 26617 34085 26651 34119
rect 27813 34085 27847 34119
rect 30297 34085 30331 34119
rect 26801 34017 26835 34051
rect 27905 34017 27939 34051
rect 28457 34017 28491 34051
rect 24593 33949 24627 33983
rect 24777 33949 24811 33983
rect 26525 33949 26559 33983
rect 27629 33949 27663 33983
rect 27721 33949 27755 33983
rect 28365 33949 28399 33983
rect 28549 33949 28583 33983
rect 29009 33949 29043 33983
rect 29193 33949 29227 33983
rect 30573 33949 30607 33983
rect 31033 33949 31067 33983
rect 31217 33949 31251 33983
rect 30297 33881 30331 33915
rect 31125 33881 31159 33915
rect 24685 33813 24719 33847
rect 26801 33813 26835 33847
rect 29101 33813 29135 33847
rect 30481 33813 30515 33847
rect 24225 33609 24259 33643
rect 26525 33609 26559 33643
rect 31233 33609 31267 33643
rect 29285 33541 29319 33575
rect 31033 33541 31067 33575
rect 23857 33473 23891 33507
rect 24869 33473 24903 33507
rect 26157 33473 26191 33507
rect 27353 33473 27387 33507
rect 27629 33473 27663 33507
rect 28365 33473 28399 33507
rect 30113 33473 30147 33507
rect 30481 33473 30515 33507
rect 30573 33473 30607 33507
rect 23949 33405 23983 33439
rect 24685 33405 24719 33439
rect 26065 33405 26099 33439
rect 27445 33405 27479 33439
rect 28457 33405 28491 33439
rect 30297 33405 30331 33439
rect 33517 33405 33551 33439
rect 25053 33337 25087 33371
rect 27169 33337 27203 33371
rect 27537 33337 27571 33371
rect 28733 33337 28767 33371
rect 33885 33337 33919 33371
rect 29377 33269 29411 33303
rect 31217 33269 31251 33303
rect 31401 33269 31435 33303
rect 33977 33269 34011 33303
rect 26709 33065 26743 33099
rect 27721 33065 27755 33099
rect 29193 33065 29227 33099
rect 30757 33065 30791 33099
rect 31309 33065 31343 33099
rect 33977 33065 34011 33099
rect 23765 32997 23799 33031
rect 25237 32997 25271 33031
rect 35173 32997 35207 33031
rect 23305 32929 23339 32963
rect 26525 32929 26559 32963
rect 27813 32929 27847 32963
rect 31493 32929 31527 32963
rect 33517 32929 33551 32963
rect 34069 32929 34103 32963
rect 35357 32929 35391 32963
rect 23029 32861 23063 32895
rect 23121 32861 23155 32895
rect 23765 32861 23799 32895
rect 24041 32861 24075 32895
rect 25145 32861 25179 32895
rect 25329 32861 25363 32895
rect 25421 32861 25455 32895
rect 26985 32861 27019 32895
rect 27537 32861 27571 32895
rect 27629 32861 27663 32895
rect 28825 32861 28859 32895
rect 31217 32861 31251 32895
rect 33701 32861 33735 32895
rect 33793 32861 33827 32895
rect 23305 32793 23339 32827
rect 29009 32793 29043 32827
rect 30389 32793 30423 32827
rect 30573 32793 30607 32827
rect 34897 32793 34931 32827
rect 23949 32725 23983 32759
rect 24961 32725 24995 32759
rect 26893 32725 26927 32759
rect 31493 32725 31527 32759
rect 25237 32521 25271 32555
rect 25973 32521 26007 32555
rect 33425 32521 33459 32555
rect 35357 32521 35391 32555
rect 23857 32385 23891 32419
rect 24869 32385 24903 32419
rect 25697 32385 25731 32419
rect 28273 32385 28307 32419
rect 28365 32385 28399 32419
rect 28457 32385 28491 32419
rect 28641 32385 28675 32419
rect 29101 32385 29135 32419
rect 29285 32385 29319 32419
rect 30573 32385 30607 32419
rect 30665 32385 30699 32419
rect 30757 32385 30791 32419
rect 30941 32385 30975 32419
rect 33609 32385 33643 32419
rect 33701 32385 33735 32419
rect 33977 32385 34011 32419
rect 34621 32385 34655 32419
rect 35265 32385 35299 32419
rect 35449 32385 35483 32419
rect 37657 32385 37691 32419
rect 23765 32317 23799 32351
rect 24961 32317 24995 32351
rect 25973 32317 26007 32351
rect 29193 32317 29227 32351
rect 34437 32317 34471 32351
rect 24225 32249 24259 32283
rect 33885 32249 33919 32283
rect 34805 32249 34839 32283
rect 25789 32181 25823 32215
rect 27997 32181 28031 32215
rect 30297 32181 30331 32215
rect 37473 32181 37507 32215
rect 21649 31977 21683 32011
rect 32045 31977 32079 32011
rect 33885 31977 33919 32011
rect 36277 31977 36311 32011
rect 23489 31909 23523 31943
rect 27445 31909 27479 31943
rect 38117 31909 38151 31943
rect 21281 31841 21315 31875
rect 22109 31841 22143 31875
rect 24593 31841 24627 31875
rect 27905 31841 27939 31875
rect 20913 31773 20947 31807
rect 21465 31773 21499 31807
rect 22376 31773 22410 31807
rect 24869 31773 24903 31807
rect 24961 31773 24995 31807
rect 25053 31773 25087 31807
rect 25237 31773 25271 31807
rect 26065 31773 26099 31807
rect 26332 31773 26366 31807
rect 28181 31773 28215 31807
rect 28273 31773 28307 31807
rect 28365 31773 28399 31807
rect 28549 31773 28583 31807
rect 29745 31773 29779 31807
rect 30665 31773 30699 31807
rect 30921 31773 30955 31807
rect 32505 31773 32539 31807
rect 34897 31773 34931 31807
rect 36921 31773 36955 31807
rect 37657 31773 37691 31807
rect 38301 31773 38335 31807
rect 32750 31705 32784 31739
rect 35142 31705 35176 31739
rect 29929 31637 29963 31671
rect 36737 31637 36771 31671
rect 37473 31637 37507 31671
rect 31033 31433 31067 31467
rect 32413 31433 32447 31467
rect 37841 31433 37875 31467
rect 28080 31365 28114 31399
rect 33425 31365 33459 31399
rect 35808 31365 35842 31399
rect 19800 31297 19834 31331
rect 22201 31297 22235 31331
rect 27813 31297 27847 31331
rect 29653 31297 29687 31331
rect 29909 31297 29943 31331
rect 31677 31297 31711 31331
rect 32597 31297 32631 31331
rect 33241 31297 33275 31331
rect 35541 31297 35575 31331
rect 37657 31297 37691 31331
rect 19533 31229 19567 31263
rect 22477 31229 22511 31263
rect 33057 31229 33091 31263
rect 37473 31229 37507 31263
rect 20913 31093 20947 31127
rect 22017 31093 22051 31127
rect 22385 31093 22419 31127
rect 29193 31093 29227 31127
rect 31493 31093 31527 31127
rect 36921 31093 36955 31127
rect 17325 30889 17359 30923
rect 22845 30889 22879 30923
rect 25605 30889 25639 30923
rect 29745 30889 29779 30923
rect 30113 30889 30147 30923
rect 36369 30889 36403 30923
rect 25697 30821 25731 30855
rect 25789 30753 25823 30787
rect 28989 30753 29023 30787
rect 36921 30753 36955 30787
rect 1593 30685 1627 30719
rect 17049 30685 17083 30719
rect 19441 30685 19475 30719
rect 19625 30685 19659 30719
rect 20269 30685 20303 30719
rect 21465 30685 21499 30719
rect 24593 30685 24627 30719
rect 24777 30685 24811 30719
rect 25513 30685 25547 30719
rect 26249 30685 26283 30719
rect 26433 30685 26467 30719
rect 26893 30685 26927 30719
rect 27077 30685 27111 30719
rect 29193 30685 29227 30719
rect 29929 30685 29963 30719
rect 30205 30685 30239 30719
rect 31033 30685 31067 30719
rect 32873 30685 32907 30719
rect 35541 30685 35575 30719
rect 36001 30685 36035 30719
rect 36185 30685 36219 30719
rect 37188 30685 37222 30719
rect 21732 30617 21766 30651
rect 26341 30617 26375 30651
rect 28917 30617 28951 30651
rect 31300 30617 31334 30651
rect 33140 30617 33174 30651
rect 1777 30549 1811 30583
rect 17509 30549 17543 30583
rect 19809 30549 19843 30583
rect 20361 30549 20395 30583
rect 24685 30549 24719 30583
rect 27077 30549 27111 30583
rect 29101 30549 29135 30583
rect 32413 30549 32447 30583
rect 34253 30549 34287 30583
rect 35357 30549 35391 30583
rect 38301 30549 38335 30583
rect 29009 30345 29043 30379
rect 33977 30345 34011 30379
rect 36737 30345 36771 30379
rect 37841 30345 37875 30379
rect 20054 30277 20088 30311
rect 34345 30277 34379 30311
rect 35624 30277 35658 30311
rect 37657 30277 37691 30311
rect 16957 30209 16991 30243
rect 17141 30209 17175 30243
rect 17785 30209 17819 30243
rect 18613 30209 18647 30243
rect 18797 30209 18831 30243
rect 19165 30209 19199 30243
rect 19809 30209 19843 30243
rect 22477 30209 22511 30243
rect 22845 30209 22879 30243
rect 23581 30209 23615 30243
rect 23848 30209 23882 30243
rect 25605 30209 25639 30243
rect 26433 30209 26467 30243
rect 26617 30209 26651 30243
rect 27169 30209 27203 30243
rect 27436 30209 27470 30243
rect 29377 30209 29411 30243
rect 34161 30209 34195 30243
rect 34253 30209 34287 30243
rect 34483 30209 34517 30243
rect 35357 30209 35391 30243
rect 37749 30209 37783 30243
rect 17693 30141 17727 30175
rect 18889 30141 18923 30175
rect 18981 30141 19015 30175
rect 22017 30141 22051 30175
rect 22201 30141 22235 30175
rect 25513 30141 25547 30175
rect 26525 30141 26559 30175
rect 29469 30141 29503 30175
rect 34621 30141 34655 30175
rect 38025 30141 38059 30175
rect 22109 30073 22143 30107
rect 25973 30073 26007 30107
rect 28549 30073 28583 30107
rect 37473 30073 37507 30107
rect 16957 30005 16991 30039
rect 18061 30005 18095 30039
rect 19349 30005 19383 30039
rect 21189 30005 21223 30039
rect 24961 30005 24995 30039
rect 29653 30005 29687 30039
rect 16497 29801 16531 29835
rect 18797 29801 18831 29835
rect 19441 29801 19475 29835
rect 22477 29801 22511 29835
rect 22937 29801 22971 29835
rect 24869 29801 24903 29835
rect 24961 29801 24995 29835
rect 25881 29801 25915 29835
rect 26065 29801 26099 29835
rect 26709 29801 26743 29835
rect 30205 29801 30239 29835
rect 34345 29801 34379 29835
rect 35265 29801 35299 29835
rect 36277 29801 36311 29835
rect 38301 29801 38335 29835
rect 18705 29733 18739 29767
rect 17325 29665 17359 29699
rect 18889 29665 18923 29699
rect 21189 29665 21223 29699
rect 22017 29665 22051 29699
rect 22109 29665 22143 29699
rect 24961 29665 24995 29699
rect 28733 29665 28767 29699
rect 29837 29665 29871 29699
rect 36185 29665 36219 29699
rect 36921 29665 36955 29699
rect 16405 29597 16439 29631
rect 16589 29597 16623 29631
rect 17233 29597 17267 29631
rect 18613 29597 18647 29631
rect 19717 29597 19751 29631
rect 19809 29597 19843 29631
rect 19901 29597 19935 29631
rect 20085 29597 20119 29631
rect 21097 29597 21131 29631
rect 21741 29597 21775 29631
rect 21925 29597 21959 29631
rect 22293 29597 22327 29631
rect 23121 29597 23155 29631
rect 23213 29597 23247 29631
rect 24593 29597 24627 29631
rect 25605 29597 25639 29631
rect 26985 29597 27019 29631
rect 27077 29597 27111 29631
rect 27169 29597 27203 29631
rect 27353 29597 27387 29631
rect 28457 29597 28491 29631
rect 28641 29597 28675 29631
rect 28825 29597 28859 29631
rect 29009 29597 29043 29631
rect 29929 29597 29963 29631
rect 31861 29597 31895 29631
rect 31953 29597 31987 29631
rect 33977 29597 34011 29631
rect 34069 29597 34103 29631
rect 34897 29597 34931 29631
rect 36277 29597 36311 29631
rect 37188 29597 37222 29631
rect 22937 29529 22971 29563
rect 24685 29529 24719 29563
rect 33793 29529 33827 29563
rect 35081 29529 35115 29563
rect 36001 29529 36035 29563
rect 17601 29461 17635 29495
rect 29193 29461 29227 29495
rect 32137 29461 32171 29495
rect 34161 29461 34195 29495
rect 36461 29461 36495 29495
rect 16957 29257 16991 29291
rect 18889 29257 18923 29291
rect 28917 29257 28951 29291
rect 30941 29257 30975 29291
rect 34253 29257 34287 29291
rect 35633 29257 35667 29291
rect 37841 29257 37875 29291
rect 22293 29189 22327 29223
rect 23090 29189 23124 29223
rect 25881 29189 25915 29223
rect 33793 29189 33827 29223
rect 17141 29121 17175 29155
rect 17417 29121 17451 29155
rect 18705 29121 18739 29155
rect 18889 29121 18923 29155
rect 22201 29121 22235 29155
rect 22385 29121 22419 29155
rect 25697 29121 25731 29155
rect 25973 29121 26007 29155
rect 26433 29121 26467 29155
rect 26525 29121 26559 29155
rect 27997 29121 28031 29155
rect 28089 29121 28123 29155
rect 28365 29121 28399 29155
rect 28825 29121 28859 29155
rect 29009 29121 29043 29155
rect 29561 29121 29595 29155
rect 29817 29121 29851 29155
rect 31769 29121 31803 29155
rect 32781 29121 32815 29155
rect 32873 29121 32907 29155
rect 34069 29121 34103 29155
rect 35357 29121 35391 29155
rect 35449 29121 35483 29155
rect 36369 29121 36403 29155
rect 36553 29121 36587 29155
rect 37565 29121 37599 29155
rect 37657 29121 37691 29155
rect 22845 29053 22879 29087
rect 33977 29053 34011 29087
rect 17325 28985 17359 29019
rect 28273 28985 28307 29019
rect 33057 28985 33091 29019
rect 24225 28917 24259 28951
rect 25697 28917 25731 28951
rect 27813 28917 27847 28951
rect 31585 28917 31619 28951
rect 33977 28917 34011 28951
rect 36737 28917 36771 28951
rect 22293 28713 22327 28747
rect 22937 28713 22971 28747
rect 23121 28713 23155 28747
rect 23765 28713 23799 28747
rect 26433 28713 26467 28747
rect 30757 28713 30791 28747
rect 30941 28713 30975 28747
rect 32781 28713 32815 28747
rect 38117 28713 38151 28747
rect 23857 28577 23891 28611
rect 33885 28577 33919 28611
rect 19809 28509 19843 28543
rect 21649 28509 21683 28543
rect 21797 28509 21831 28543
rect 22025 28509 22059 28543
rect 22155 28509 22189 28543
rect 23581 28509 23615 28543
rect 23673 28509 23707 28543
rect 25053 28509 25087 28543
rect 27261 28509 27295 28543
rect 27537 28509 27571 28543
rect 28181 28509 28215 28543
rect 28457 28509 28491 28543
rect 28641 28509 28675 28543
rect 29929 28509 29963 28543
rect 31401 28509 31435 28543
rect 31668 28509 31702 28543
rect 33425 28509 33459 28543
rect 34069 28509 34103 28543
rect 34897 28509 34931 28543
rect 36737 28509 36771 28543
rect 20076 28441 20110 28475
rect 21925 28441 21959 28475
rect 22753 28441 22787 28475
rect 22969 28441 23003 28475
rect 25320 28441 25354 28475
rect 27445 28441 27479 28475
rect 30573 28441 30607 28475
rect 35142 28441 35176 28475
rect 36982 28441 37016 28475
rect 21189 28373 21223 28407
rect 27077 28373 27111 28407
rect 27997 28373 28031 28407
rect 30021 28373 30055 28407
rect 30773 28373 30807 28407
rect 33241 28373 33275 28407
rect 34253 28373 34287 28407
rect 36277 28373 36311 28407
rect 23581 28169 23615 28203
rect 25789 28169 25823 28203
rect 26157 28169 26191 28203
rect 27261 28169 27295 28203
rect 28641 28169 28675 28203
rect 30573 28169 30607 28203
rect 31493 28169 31527 28203
rect 33701 28169 33735 28203
rect 34805 28169 34839 28203
rect 36001 28169 36035 28203
rect 20177 28101 20211 28135
rect 28365 28101 28399 28135
rect 30297 28101 30331 28135
rect 32588 28101 32622 28135
rect 17141 28033 17175 28067
rect 18521 28033 18555 28067
rect 19717 28033 19751 28067
rect 19809 28033 19843 28067
rect 20637 28033 20671 28067
rect 20821 28033 20855 28067
rect 21281 28033 21315 28067
rect 22477 28033 22511 28067
rect 23397 28033 23431 28067
rect 24593 28033 24627 28067
rect 25973 28033 26007 28067
rect 26249 28033 26283 28067
rect 27169 28033 27203 28067
rect 27997 28033 28031 28067
rect 28090 28033 28124 28067
rect 28273 28033 28307 28067
rect 28462 28033 28496 28067
rect 29929 28033 29963 28067
rect 30022 28033 30056 28067
rect 30205 28033 30239 28067
rect 30394 28033 30428 28067
rect 31033 28033 31067 28067
rect 34345 28033 34379 28067
rect 34989 28033 35023 28067
rect 36185 28033 36219 28067
rect 36829 28033 36863 28067
rect 37657 28033 37691 28067
rect 17233 27965 17267 27999
rect 18429 27965 18463 27999
rect 20085 27965 20119 27999
rect 22753 27965 22787 27999
rect 23213 27965 23247 27999
rect 24409 27965 24443 27999
rect 32321 27965 32355 27999
rect 37473 27965 37507 27999
rect 17509 27897 17543 27931
rect 18889 27897 18923 27931
rect 19993 27897 20027 27931
rect 20637 27897 20671 27931
rect 21373 27897 21407 27931
rect 24777 27897 24811 27931
rect 34161 27897 34195 27931
rect 22293 27829 22327 27863
rect 22661 27829 22695 27863
rect 31125 27829 31159 27863
rect 36645 27829 36679 27863
rect 37841 27829 37875 27863
rect 18337 27625 18371 27659
rect 23121 27625 23155 27659
rect 27077 27625 27111 27659
rect 34345 27625 34379 27659
rect 35633 27625 35667 27659
rect 16865 27557 16899 27591
rect 17325 27557 17359 27591
rect 17693 27557 17727 27591
rect 23581 27557 23615 27591
rect 25697 27557 25731 27591
rect 30481 27557 30515 27591
rect 33425 27557 33459 27591
rect 16589 27489 16623 27523
rect 17601 27489 17635 27523
rect 27813 27489 27847 27523
rect 30113 27489 30147 27523
rect 36645 27489 36679 27523
rect 16497 27421 16531 27455
rect 17509 27421 17543 27455
rect 17785 27421 17819 27455
rect 18613 27421 18647 27455
rect 21741 27421 21775 27455
rect 22008 27421 22042 27455
rect 23581 27421 23615 27455
rect 23765 27421 23799 27455
rect 24593 27421 24627 27455
rect 24777 27421 24811 27455
rect 25973 27421 26007 27455
rect 26525 27421 26559 27455
rect 26801 27421 26835 27455
rect 26893 27421 26927 27455
rect 27537 27421 27571 27455
rect 27721 27421 27755 27455
rect 27905 27421 27939 27455
rect 28089 27421 28123 27455
rect 29193 27421 29227 27455
rect 29745 27421 29779 27455
rect 29929 27421 29963 27455
rect 30021 27421 30055 27455
rect 30297 27421 30331 27455
rect 31217 27421 31251 27455
rect 34069 27421 34103 27455
rect 34161 27421 34195 27455
rect 35081 27421 35115 27455
rect 35633 27421 35667 27455
rect 35817 27421 35851 27455
rect 36901 27421 36935 27455
rect 18337 27353 18371 27387
rect 25697 27353 25731 27387
rect 26709 27353 26743 27387
rect 31462 27353 31496 27387
rect 33149 27353 33183 27387
rect 18521 27285 18555 27319
rect 24685 27285 24719 27319
rect 25881 27285 25915 27319
rect 28273 27285 28307 27319
rect 29009 27285 29043 27319
rect 32597 27285 32631 27319
rect 34897 27285 34931 27319
rect 36001 27285 36035 27319
rect 38025 27285 38059 27319
rect 17325 27081 17359 27115
rect 22753 27081 22787 27115
rect 25329 27081 25363 27115
rect 26357 27081 26391 27115
rect 27261 27081 27295 27115
rect 28825 27081 28859 27115
rect 30481 27081 30515 27115
rect 32597 27081 32631 27115
rect 33885 27081 33919 27115
rect 35725 27081 35759 27115
rect 37841 27081 37875 27115
rect 18613 27013 18647 27047
rect 19962 27013 19996 27047
rect 24216 27013 24250 27047
rect 26157 27013 26191 27047
rect 28457 27013 28491 27047
rect 31585 27013 31619 27047
rect 31769 27013 31803 27047
rect 17049 26945 17083 26979
rect 17969 26945 18003 26979
rect 18889 26945 18923 26979
rect 18981 26945 19015 26979
rect 19073 26945 19107 26979
rect 19257 26945 19291 26979
rect 22017 26945 22051 26979
rect 22201 26945 22235 26979
rect 22569 26945 22603 26979
rect 27169 26945 27203 26979
rect 28181 26945 28215 26979
rect 28274 26945 28308 26979
rect 28549 26945 28583 26979
rect 28687 26945 28721 26979
rect 29561 26945 29595 26979
rect 30297 26945 30331 26979
rect 30573 26945 30607 26979
rect 32505 26945 32539 26979
rect 33701 26945 33735 26979
rect 34345 26945 34379 26979
rect 34612 26945 34646 26979
rect 36369 26945 36403 26979
rect 36461 26945 36495 26979
rect 36645 26945 36679 26979
rect 37473 26945 37507 26979
rect 37657 26945 37691 26979
rect 17325 26877 17359 26911
rect 17785 26877 17819 26911
rect 19717 26877 19751 26911
rect 22293 26877 22327 26911
rect 22385 26877 22419 26911
rect 23949 26877 23983 26911
rect 29837 26877 29871 26911
rect 33517 26877 33551 26911
rect 17141 26809 17175 26843
rect 36553 26809 36587 26843
rect 18153 26741 18187 26775
rect 21097 26741 21131 26775
rect 26341 26741 26375 26775
rect 26525 26741 26559 26775
rect 30297 26741 30331 26775
rect 36185 26741 36219 26775
rect 17877 26537 17911 26571
rect 18613 26537 18647 26571
rect 18705 26537 18739 26571
rect 21373 26537 21407 26571
rect 26525 26537 26559 26571
rect 27445 26537 27479 26571
rect 28089 26537 28123 26571
rect 29009 26537 29043 26571
rect 36277 26537 36311 26571
rect 36461 26469 36495 26503
rect 38301 26469 38335 26503
rect 18797 26401 18831 26435
rect 30389 26401 30423 26435
rect 33425 26401 33459 26435
rect 35541 26401 35575 26435
rect 36921 26401 36955 26435
rect 17877 26333 17911 26367
rect 18061 26333 18095 26367
rect 18521 26333 18555 26367
rect 21281 26333 21315 26367
rect 22937 26333 22971 26367
rect 23121 26333 23155 26367
rect 25145 26333 25179 26367
rect 27353 26333 27387 26367
rect 27997 26333 28031 26367
rect 28917 26333 28951 26367
rect 30113 26333 30147 26367
rect 30297 26333 30331 26367
rect 33609 26333 33643 26367
rect 35081 26333 35115 26367
rect 35173 26333 35207 26367
rect 35265 26333 35299 26367
rect 25412 26265 25446 26299
rect 29929 26265 29963 26299
rect 31217 26265 31251 26299
rect 33793 26265 33827 26299
rect 35383 26265 35417 26299
rect 36093 26265 36127 26299
rect 37166 26265 37200 26299
rect 23029 26197 23063 26231
rect 32505 26197 32539 26231
rect 34897 26197 34931 26231
rect 36303 26197 36337 26231
rect 22937 25993 22971 26027
rect 24685 25993 24719 26027
rect 25605 25993 25639 26027
rect 34345 25993 34379 26027
rect 36093 25993 36127 26027
rect 22569 25925 22603 25959
rect 22785 25925 22819 25959
rect 30104 25925 30138 25959
rect 32413 25925 32447 25959
rect 37841 25925 37875 25959
rect 17601 25857 17635 25891
rect 19717 25857 19751 25891
rect 19809 25857 19843 25891
rect 19901 25857 19935 25891
rect 20085 25857 20119 25891
rect 23397 25857 23431 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 29101 25857 29135 25891
rect 32321 25857 32355 25891
rect 32965 25857 32999 25891
rect 33232 25857 33266 25891
rect 34989 25857 35023 25891
rect 36277 25857 36311 25891
rect 36921 25857 36955 25891
rect 37657 25857 37691 25891
rect 17509 25789 17543 25823
rect 25881 25789 25915 25823
rect 29377 25789 29411 25823
rect 29837 25789 29871 25823
rect 34805 25789 34839 25823
rect 37473 25789 37507 25823
rect 17969 25721 18003 25755
rect 31217 25721 31251 25755
rect 19441 25653 19475 25687
rect 22753 25653 22787 25687
rect 29193 25653 29227 25687
rect 29285 25653 29319 25687
rect 35173 25653 35207 25687
rect 36737 25653 36771 25687
rect 17233 25449 17267 25483
rect 21189 25449 21223 25483
rect 22201 25449 22235 25483
rect 25513 25449 25547 25483
rect 27169 25449 27203 25483
rect 29009 25449 29043 25483
rect 31401 25449 31435 25483
rect 34069 25449 34103 25483
rect 24041 25381 24075 25415
rect 24777 25381 24811 25415
rect 27353 25381 27387 25415
rect 17509 25313 17543 25347
rect 17601 25313 17635 25347
rect 18613 25313 18647 25347
rect 24869 25313 24903 25347
rect 25605 25313 25639 25347
rect 26157 25313 26191 25347
rect 30021 25313 30055 25347
rect 36921 25313 36955 25347
rect 17417 25245 17451 25279
rect 17693 25245 17727 25279
rect 18245 25245 18279 25279
rect 18705 25245 18739 25279
rect 19809 25245 19843 25279
rect 20076 25245 20110 25279
rect 21649 25245 21683 25279
rect 21833 25245 21867 25279
rect 22017 25245 22051 25279
rect 22661 25245 22695 25279
rect 22928 25245 22962 25279
rect 24593 25245 24627 25279
rect 24685 25245 24719 25279
rect 25329 25245 25363 25279
rect 25421 25245 25455 25279
rect 26341 25245 26375 25279
rect 27813 25245 27847 25279
rect 27997 25245 28031 25279
rect 32045 25245 32079 25279
rect 33885 25245 33919 25279
rect 34897 25245 34931 25279
rect 37177 25245 37211 25279
rect 21925 25177 21959 25211
rect 26985 25177 27019 25211
rect 28825 25177 28859 25211
rect 29041 25177 29075 25211
rect 30288 25177 30322 25211
rect 32312 25177 32346 25211
rect 35142 25177 35176 25211
rect 18889 25109 18923 25143
rect 26525 25109 26559 25143
rect 27185 25109 27219 25143
rect 27905 25109 27939 25143
rect 29193 25109 29227 25143
rect 33425 25109 33459 25143
rect 36277 25109 36311 25143
rect 38301 25109 38335 25143
rect 24869 24905 24903 24939
rect 28549 24905 28583 24939
rect 34897 24905 34931 24939
rect 37657 24905 37691 24939
rect 22201 24837 22235 24871
rect 22937 24837 22971 24871
rect 37841 24837 37875 24871
rect 16129 24769 16163 24803
rect 16313 24769 16347 24803
rect 17049 24769 17083 24803
rect 17785 24769 17819 24803
rect 17969 24769 18003 24803
rect 18613 24769 18647 24803
rect 18889 24769 18923 24803
rect 19073 24769 19107 24803
rect 20168 24769 20202 24803
rect 22017 24769 22051 24803
rect 22845 24769 22879 24803
rect 23489 24769 23523 24803
rect 23756 24769 23790 24803
rect 25329 24769 25363 24803
rect 25513 24769 25547 24803
rect 25973 24769 26007 24803
rect 27169 24769 27203 24803
rect 27436 24769 27470 24803
rect 29265 24769 29299 24803
rect 30849 24769 30883 24803
rect 31033 24769 31067 24803
rect 31677 24769 31711 24803
rect 32597 24769 32631 24803
rect 32873 24769 32907 24803
rect 33701 24769 33735 24803
rect 35081 24769 35115 24803
rect 36461 24769 36495 24803
rect 36737 24769 36771 24803
rect 37473 24769 37507 24803
rect 37749 24769 37783 24803
rect 16221 24701 16255 24735
rect 17325 24701 17359 24735
rect 19901 24701 19935 24735
rect 22385 24701 22419 24735
rect 26249 24701 26283 24735
rect 29009 24701 29043 24735
rect 32781 24701 32815 24735
rect 36645 24701 36679 24735
rect 17233 24633 17267 24667
rect 18889 24633 18923 24667
rect 26157 24633 26191 24667
rect 30849 24633 30883 24667
rect 33517 24633 33551 24667
rect 36921 24633 36955 24667
rect 38025 24633 38059 24667
rect 17141 24565 17175 24599
rect 18153 24565 18187 24599
rect 21281 24565 21315 24599
rect 25329 24565 25363 24599
rect 26065 24565 26099 24599
rect 30389 24565 30423 24599
rect 31493 24565 31527 24599
rect 32597 24565 32631 24599
rect 33057 24565 33091 24599
rect 36737 24565 36771 24599
rect 17049 24361 17083 24395
rect 17141 24361 17175 24395
rect 19533 24361 19567 24395
rect 22293 24361 22327 24395
rect 24593 24361 24627 24395
rect 27261 24361 27295 24395
rect 27353 24361 27387 24395
rect 28549 24361 28583 24395
rect 28917 24361 28951 24395
rect 30113 24361 30147 24395
rect 33425 24361 33459 24395
rect 37565 24361 37599 24395
rect 18797 24293 18831 24327
rect 23765 24293 23799 24327
rect 26709 24293 26743 24327
rect 17233 24225 17267 24259
rect 17969 24225 18003 24259
rect 21097 24225 21131 24259
rect 22937 24225 22971 24259
rect 25329 24225 25363 24259
rect 27445 24225 27479 24259
rect 33885 24225 33919 24259
rect 36185 24225 36219 24259
rect 16957 24157 16991 24191
rect 17877 24157 17911 24191
rect 18705 24157 18739 24191
rect 18889 24157 18923 24191
rect 19809 24157 19843 24191
rect 19901 24157 19935 24191
rect 19993 24157 20027 24191
rect 20177 24157 20211 24191
rect 21005 24157 21039 24191
rect 21649 24157 21683 24191
rect 21742 24157 21776 24191
rect 22017 24157 22051 24191
rect 22155 24157 22189 24191
rect 23121 24157 23155 24191
rect 23305 24157 23339 24191
rect 24041 24157 24075 24191
rect 24593 24157 24627 24191
rect 24777 24157 24811 24191
rect 25585 24157 25619 24191
rect 27169 24157 27203 24191
rect 28733 24157 28767 24191
rect 29009 24157 29043 24191
rect 29745 24157 29779 24191
rect 29929 24157 29963 24191
rect 30665 24157 30699 24191
rect 30757 24157 30791 24191
rect 30941 24157 30975 24191
rect 31585 24157 31619 24191
rect 32045 24157 32079 24191
rect 32301 24157 32335 24191
rect 34069 24157 34103 24191
rect 34253 24157 34287 24191
rect 35081 24157 35115 24191
rect 21925 24089 21959 24123
rect 23765 24089 23799 24123
rect 36452 24089 36486 24123
rect 18245 24021 18279 24055
rect 23949 24021 23983 24055
rect 31401 24021 31435 24055
rect 34897 24021 34931 24055
rect 17969 23817 18003 23851
rect 19441 23817 19475 23851
rect 22753 23817 22787 23851
rect 29101 23817 29135 23851
rect 36645 23817 36679 23851
rect 17877 23749 17911 23783
rect 23397 23749 23431 23783
rect 30472 23749 30506 23783
rect 35541 23749 35575 23783
rect 19257 23681 19291 23715
rect 19441 23681 19475 23715
rect 21281 23681 21315 23715
rect 22017 23681 22051 23715
rect 22201 23681 22235 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 25973 23681 26007 23715
rect 26065 23681 26099 23715
rect 26341 23681 26375 23715
rect 29009 23681 29043 23715
rect 29193 23681 29227 23715
rect 32873 23681 32907 23715
rect 33057 23681 33091 23715
rect 33793 23681 33827 23715
rect 36829 23681 36863 23715
rect 37473 23681 37507 23715
rect 37657 23681 37691 23715
rect 22293 23613 22327 23647
rect 25789 23613 25823 23647
rect 30205 23613 30239 23647
rect 32781 23613 32815 23647
rect 32965 23613 32999 23647
rect 24685 23545 24719 23579
rect 21373 23477 21407 23511
rect 26249 23477 26283 23511
rect 31585 23477 31619 23511
rect 32597 23477 32631 23511
rect 37841 23477 37875 23511
rect 19625 23273 19659 23307
rect 21373 23273 21407 23307
rect 24041 23273 24075 23307
rect 25881 23273 25915 23307
rect 29009 23273 29043 23307
rect 31217 23273 31251 23307
rect 34069 23273 34103 23307
rect 34253 23273 34287 23307
rect 38301 23273 38335 23307
rect 32321 23205 32355 23239
rect 32781 23205 32815 23239
rect 20821 23137 20855 23171
rect 22661 23137 22695 23171
rect 25329 23137 25363 23171
rect 26341 23137 26375 23171
rect 31953 23137 31987 23171
rect 36921 23137 36955 23171
rect 17785 23069 17819 23103
rect 17969 23069 18003 23103
rect 19441 23069 19475 23103
rect 20729 23069 20763 23103
rect 21557 23069 21591 23103
rect 21649 23069 21683 23103
rect 21833 23069 21867 23103
rect 21935 23069 21969 23103
rect 25053 23069 25087 23103
rect 25145 23069 25179 23103
rect 26065 23069 26099 23103
rect 26157 23069 26191 23103
rect 26433 23069 26467 23103
rect 26893 23069 26927 23103
rect 27077 23069 27111 23103
rect 27629 23069 27663 23103
rect 32137 23069 32171 23103
rect 33057 23069 33091 23103
rect 33149 23069 33183 23103
rect 33246 23069 33280 23103
rect 33425 23069 33459 23103
rect 34897 23069 34931 23103
rect 18429 23001 18463 23035
rect 18613 23001 18647 23035
rect 22928 23001 22962 23035
rect 26985 23001 27019 23035
rect 27896 23001 27930 23035
rect 29745 23001 29779 23035
rect 33885 23001 33919 23035
rect 35142 23001 35176 23035
rect 37188 23001 37222 23035
rect 17969 22933 18003 22967
rect 18797 22933 18831 22967
rect 34095 22933 34129 22967
rect 36277 22933 36311 22967
rect 17877 22729 17911 22763
rect 17969 22729 18003 22763
rect 21005 22729 21039 22763
rect 23397 22729 23431 22763
rect 25697 22729 25731 22763
rect 26617 22729 26651 22763
rect 30573 22729 30607 22763
rect 33701 22729 33735 22763
rect 34253 22729 34287 22763
rect 37841 22729 37875 22763
rect 19870 22661 19904 22695
rect 22569 22661 22603 22695
rect 22785 22661 22819 22695
rect 23673 22661 23707 22695
rect 32588 22661 32622 22695
rect 35142 22661 35176 22695
rect 17601 22593 17635 22627
rect 18061 22593 18095 22627
rect 18797 22593 18831 22627
rect 18886 22599 18920 22633
rect 18981 22596 19015 22630
rect 19165 22593 19199 22627
rect 23397 22593 23431 22627
rect 23489 22593 23523 22627
rect 24584 22593 24618 22627
rect 27988 22593 28022 22627
rect 29745 22593 29779 22627
rect 30297 22593 30331 22627
rect 31309 22593 31343 22627
rect 32321 22593 32355 22627
rect 34437 22593 34471 22627
rect 34897 22593 34931 22627
rect 37565 22593 37599 22627
rect 37657 22593 37691 22627
rect 19625 22525 19659 22559
rect 24317 22525 24351 22559
rect 26157 22525 26191 22559
rect 27721 22525 27755 22559
rect 31125 22525 31159 22559
rect 18521 22457 18555 22491
rect 22937 22457 22971 22491
rect 26433 22457 26467 22491
rect 29101 22457 29135 22491
rect 29561 22457 29595 22491
rect 22753 22389 22787 22423
rect 31493 22389 31527 22423
rect 36277 22389 36311 22423
rect 18613 22185 18647 22219
rect 20453 22185 20487 22219
rect 22477 22185 22511 22219
rect 24777 22185 24811 22219
rect 29009 22185 29043 22219
rect 33333 22185 33367 22219
rect 34345 22185 34379 22219
rect 36001 22185 36035 22219
rect 37381 22185 37415 22219
rect 21005 22117 21039 22151
rect 23029 22117 23063 22151
rect 26893 22117 26927 22151
rect 26985 22117 27019 22151
rect 28365 22117 28399 22151
rect 17765 22049 17799 22083
rect 26065 22049 26099 22083
rect 26525 22049 26559 22083
rect 32413 22049 32447 22083
rect 34989 22049 35023 22083
rect 35541 22049 35575 22083
rect 36185 22049 36219 22083
rect 17969 21981 18003 22015
rect 20269 21981 20303 22015
rect 20545 21981 20579 22015
rect 21189 21981 21223 22015
rect 21281 21981 21315 22015
rect 22293 21981 22327 22015
rect 22569 21981 22603 22015
rect 23305 21981 23339 22015
rect 24961 21981 24995 22015
rect 25789 21981 25823 22015
rect 25881 21981 25915 22015
rect 28549 21981 28583 22015
rect 29193 21981 29227 22015
rect 30021 21981 30055 22015
rect 32321 21981 32355 22015
rect 32505 21981 32539 22015
rect 32597 21981 32631 22015
rect 34069 21981 34103 22015
rect 34161 21981 34195 22015
rect 35265 21981 35299 22015
rect 36277 21981 36311 22015
rect 37565 21981 37599 22015
rect 17693 21913 17727 21947
rect 17877 21913 17911 21947
rect 18429 21913 18463 21947
rect 18629 21913 18663 21947
rect 21005 21913 21039 21947
rect 23029 21913 23063 21947
rect 30288 21913 30322 21947
rect 33241 21913 33275 21947
rect 35173 21913 35207 21947
rect 36001 21913 36035 21947
rect 18797 21845 18831 21879
rect 20085 21845 20119 21879
rect 22109 21845 22143 21879
rect 23213 21845 23247 21879
rect 31401 21845 31435 21879
rect 32137 21845 32171 21879
rect 35357 21845 35391 21879
rect 36461 21845 36495 21879
rect 18889 21641 18923 21675
rect 21189 21641 21223 21675
rect 23397 21641 23431 21675
rect 27997 21641 28031 21675
rect 29377 21641 29411 21675
rect 32321 21641 32355 21675
rect 33609 21641 33643 21675
rect 36645 21641 36679 21675
rect 22262 21573 22296 21607
rect 27537 21573 27571 21607
rect 30113 21573 30147 21607
rect 31033 21573 31067 21607
rect 33517 21573 33551 21607
rect 34805 21573 34839 21607
rect 18613 21505 18647 21539
rect 18705 21505 18739 21539
rect 19809 21505 19843 21539
rect 20076 21505 20110 21539
rect 22017 21505 22051 21539
rect 23857 21505 23891 21539
rect 24041 21505 24075 21539
rect 24777 21505 24811 21539
rect 25881 21505 25915 21539
rect 26617 21505 26651 21539
rect 27353 21505 27387 21539
rect 28273 21505 28307 21539
rect 29193 21505 29227 21539
rect 32597 21505 32631 21539
rect 32689 21505 32723 21539
rect 32781 21505 32815 21539
rect 32965 21505 32999 21539
rect 34529 21505 34563 21539
rect 34621 21505 34655 21539
rect 35532 21505 35566 21539
rect 18889 21437 18923 21471
rect 27169 21437 27203 21471
rect 28181 21437 28215 21471
rect 28365 21437 28399 21471
rect 28457 21437 28491 21471
rect 29009 21437 29043 21471
rect 35265 21437 35299 21471
rect 30389 21369 30423 21403
rect 23857 21301 23891 21335
rect 25053 21301 25087 21335
rect 25697 21301 25731 21335
rect 26433 21301 26467 21335
rect 31125 21301 31159 21335
rect 23857 21097 23891 21131
rect 28825 21097 28859 21131
rect 27813 21029 27847 21063
rect 24593 20961 24627 20995
rect 30297 20961 30331 20995
rect 1777 20893 1811 20927
rect 22477 20893 22511 20927
rect 26433 20893 26467 20927
rect 28641 20893 28675 20927
rect 30564 20893 30598 20927
rect 32689 20893 32723 20927
rect 34897 20893 34931 20927
rect 22744 20825 22778 20859
rect 24860 20825 24894 20859
rect 26700 20825 26734 20859
rect 28273 20825 28307 20859
rect 32956 20825 32990 20859
rect 35164 20825 35198 20859
rect 25973 20757 26007 20791
rect 28457 20757 28491 20791
rect 28549 20757 28583 20791
rect 31677 20757 31711 20791
rect 34069 20757 34103 20791
rect 36277 20757 36311 20791
rect 24409 20553 24443 20587
rect 31309 20553 31343 20587
rect 32781 20553 32815 20587
rect 34069 20553 34103 20587
rect 36001 20553 36035 20587
rect 36645 20553 36679 20587
rect 19717 20485 19751 20519
rect 29000 20485 29034 20519
rect 32321 20485 32355 20519
rect 35541 20485 35575 20519
rect 20545 20417 20579 20451
rect 20729 20417 20763 20451
rect 24317 20417 24351 20451
rect 24501 20417 24535 20451
rect 25237 20417 25271 20451
rect 25504 20417 25538 20451
rect 27905 20417 27939 20451
rect 27997 20417 28031 20451
rect 28181 20417 28215 20451
rect 31033 20417 31067 20451
rect 31125 20417 31159 20451
rect 32597 20417 32631 20451
rect 33425 20417 33459 20451
rect 33609 20417 33643 20451
rect 34253 20417 34287 20451
rect 35265 20417 35299 20451
rect 35357 20417 35391 20451
rect 36185 20417 36219 20451
rect 36829 20417 36863 20451
rect 28733 20349 28767 20383
rect 32505 20349 32539 20383
rect 33241 20349 33275 20383
rect 26617 20281 26651 20315
rect 28089 20281 28123 20315
rect 19993 20213 20027 20247
rect 20545 20213 20579 20247
rect 27721 20213 27755 20247
rect 30113 20213 30147 20247
rect 32321 20213 32355 20247
rect 26249 20009 26283 20043
rect 28365 20009 28399 20043
rect 28641 20009 28675 20043
rect 33885 20009 33919 20043
rect 24869 19941 24903 19975
rect 25881 19873 25915 19907
rect 31125 19873 31159 19907
rect 19901 19805 19935 19839
rect 22201 19805 22235 19839
rect 22385 19805 22419 19839
rect 23857 19805 23891 19839
rect 24041 19805 24075 19839
rect 25145 19805 25179 19839
rect 26065 19805 26099 19839
rect 28273 19805 28307 19839
rect 28457 19805 28491 19839
rect 29745 19805 29779 19839
rect 29929 19805 29963 19839
rect 31309 19805 31343 19839
rect 32505 19805 32539 19839
rect 34989 19805 35023 19839
rect 35081 19805 35115 19839
rect 36001 19805 36035 19839
rect 20168 19737 20202 19771
rect 24869 19737 24903 19771
rect 32772 19737 32806 19771
rect 21281 19669 21315 19703
rect 22293 19669 22327 19703
rect 23949 19669 23983 19703
rect 25053 19669 25087 19703
rect 30113 19669 30147 19703
rect 31493 19669 31527 19703
rect 35265 19669 35299 19703
rect 35817 19669 35851 19703
rect 20361 19465 20395 19499
rect 25605 19465 25639 19499
rect 26065 19465 26099 19499
rect 28641 19465 28675 19499
rect 30757 19465 30791 19499
rect 32781 19465 32815 19499
rect 33441 19465 33475 19499
rect 33609 19465 33643 19499
rect 37473 19465 37507 19499
rect 22284 19397 22318 19431
rect 24492 19397 24526 19431
rect 31769 19397 31803 19431
rect 33241 19397 33275 19431
rect 35808 19397 35842 19431
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 20545 19329 20579 19363
rect 22017 19329 22051 19363
rect 26249 19329 26283 19363
rect 27353 19329 27387 19363
rect 28181 19329 28215 19363
rect 28457 19329 28491 19363
rect 29469 19329 29503 19363
rect 30113 19329 30147 19363
rect 30941 19329 30975 19363
rect 31585 19329 31619 19363
rect 32321 19329 32355 19363
rect 32597 19329 32631 19363
rect 34713 19329 34747 19363
rect 37657 19329 37691 19363
rect 20821 19261 20855 19295
rect 24225 19261 24259 19295
rect 28365 19261 28399 19295
rect 31401 19261 31435 19295
rect 32505 19261 32539 19295
rect 35541 19261 35575 19295
rect 19717 19125 19751 19159
rect 20729 19125 20763 19159
rect 23397 19125 23431 19159
rect 27169 19125 27203 19159
rect 28457 19125 28491 19159
rect 29285 19125 29319 19159
rect 29929 19125 29963 19159
rect 32505 19125 32539 19159
rect 33425 19125 33459 19159
rect 34529 19125 34563 19159
rect 36921 19125 36955 19159
rect 25973 18921 26007 18955
rect 28825 18921 28859 18955
rect 33425 18921 33459 18955
rect 32965 18785 32999 18819
rect 19625 18717 19659 18751
rect 19881 18717 19915 18751
rect 21465 18717 21499 18751
rect 21649 18717 21683 18751
rect 22569 18717 22603 18751
rect 24593 18717 24627 18751
rect 26433 18717 26467 18751
rect 28273 18717 28307 18751
rect 28549 18717 28583 18751
rect 31217 18717 31251 18751
rect 33609 18717 33643 18751
rect 34253 18717 34287 18751
rect 34897 18717 34931 18751
rect 36737 18717 36771 18751
rect 37004 18717 37038 18751
rect 21833 18649 21867 18683
rect 22836 18649 22870 18683
rect 24860 18649 24894 18683
rect 26700 18649 26734 18683
rect 28457 18649 28491 18683
rect 35142 18649 35176 18683
rect 21005 18581 21039 18615
rect 23949 18581 23983 18615
rect 27813 18581 27847 18615
rect 28641 18581 28675 18615
rect 34069 18581 34103 18615
rect 36277 18581 36311 18615
rect 38117 18581 38151 18615
rect 20177 18377 20211 18411
rect 20837 18377 20871 18411
rect 22661 18377 22695 18411
rect 24685 18377 24719 18411
rect 25605 18377 25639 18411
rect 28549 18377 28583 18411
rect 31125 18377 31159 18411
rect 33793 18377 33827 18411
rect 36001 18377 36035 18411
rect 20637 18309 20671 18343
rect 32680 18309 32714 18343
rect 34713 18309 34747 18343
rect 34805 18309 34839 18343
rect 37473 18309 37507 18343
rect 37673 18309 37707 18343
rect 19901 18241 19935 18275
rect 19993 18241 20027 18275
rect 22385 18241 22419 18275
rect 23397 18241 23431 18275
rect 25789 18241 25823 18275
rect 26065 18241 26099 18275
rect 27169 18241 27203 18275
rect 27425 18241 27459 18275
rect 29745 18241 29779 18275
rect 30001 18241 30035 18275
rect 32413 18241 32447 18275
rect 34621 18241 34655 18275
rect 34923 18241 34957 18275
rect 35725 18241 35759 18275
rect 35817 18241 35851 18275
rect 36461 18241 36495 18275
rect 36645 18241 36679 18275
rect 20177 18173 20211 18207
rect 22661 18173 22695 18207
rect 35081 18173 35115 18207
rect 21005 18105 21039 18139
rect 37841 18105 37875 18139
rect 20821 18037 20855 18071
rect 22477 18037 22511 18071
rect 25973 18037 26007 18071
rect 34437 18037 34471 18071
rect 36553 18037 36587 18071
rect 36829 18037 36863 18071
rect 37657 18037 37691 18071
rect 20361 17833 20395 17867
rect 22477 17833 22511 17867
rect 23489 17833 23523 17867
rect 25973 17833 26007 17867
rect 26985 17833 27019 17867
rect 29745 17833 29779 17867
rect 32505 17833 32539 17867
rect 33793 17833 33827 17867
rect 35265 17833 35299 17867
rect 36921 17833 36955 17867
rect 20913 17765 20947 17799
rect 22661 17765 22695 17799
rect 35541 17765 35575 17799
rect 26617 17697 26651 17731
rect 27445 17697 27479 17731
rect 30389 17697 30423 17731
rect 20177 17629 20211 17663
rect 20453 17629 20487 17663
rect 21189 17629 21223 17663
rect 23121 17629 23155 17663
rect 23305 17629 23339 17663
rect 24685 17629 24719 17663
rect 24778 17629 24812 17663
rect 24915 17629 24949 17663
rect 25150 17629 25184 17663
rect 26801 17629 26835 17663
rect 27629 17629 27663 17663
rect 28825 17629 28859 17663
rect 28917 17629 28951 17663
rect 29929 17629 29963 17663
rect 30573 17629 30607 17663
rect 31217 17629 31251 17663
rect 33425 17629 33459 17663
rect 33609 17629 33643 17663
rect 35449 17629 35483 17663
rect 35633 17629 35667 17663
rect 35761 17629 35795 17663
rect 36645 17629 36679 17663
rect 36737 17629 36771 17663
rect 37473 17629 37507 17663
rect 37565 17629 37599 17663
rect 20913 17561 20947 17595
rect 22293 17561 22327 17595
rect 22509 17561 22543 17595
rect 25053 17561 25087 17595
rect 25789 17561 25823 17595
rect 25989 17561 26023 17595
rect 27813 17561 27847 17595
rect 19993 17493 20027 17527
rect 21097 17493 21131 17527
rect 25329 17493 25363 17527
rect 26157 17493 26191 17527
rect 29101 17493 29135 17527
rect 30757 17493 30791 17527
rect 37749 17493 37783 17527
rect 22937 17289 22971 17323
rect 24685 17289 24719 17323
rect 26525 17289 26559 17323
rect 29745 17289 29779 17323
rect 32873 17289 32907 17323
rect 34805 17289 34839 17323
rect 36829 17289 36863 17323
rect 19800 17221 19834 17255
rect 23397 17221 23431 17255
rect 26341 17221 26375 17255
rect 27169 17221 27203 17255
rect 27353 17221 27387 17255
rect 30472 17221 30506 17255
rect 32321 17221 32355 17255
rect 32505 17221 32539 17255
rect 33692 17221 33726 17255
rect 36369 17221 36403 17255
rect 19533 17153 19567 17187
rect 22661 17153 22695 17187
rect 22753 17153 22787 17187
rect 25605 17153 25639 17187
rect 26617 17153 26651 17187
rect 27445 17153 27479 17187
rect 28365 17153 28399 17187
rect 28621 17153 28655 17187
rect 30205 17153 30239 17187
rect 32597 17153 32631 17187
rect 32689 17153 32723 17187
rect 35449 17153 35483 17187
rect 36645 17153 36679 17187
rect 37657 17153 37691 17187
rect 22937 17085 22971 17119
rect 25881 17085 25915 17119
rect 33425 17085 33459 17119
rect 36461 17085 36495 17119
rect 25697 17017 25731 17051
rect 26341 17017 26375 17051
rect 31585 17017 31619 17051
rect 20913 16949 20947 16983
rect 25605 16949 25639 16983
rect 27169 16949 27203 16983
rect 35265 16949 35299 16983
rect 36553 16949 36587 16983
rect 37473 16949 37507 16983
rect 25697 16745 25731 16779
rect 28365 16745 28399 16779
rect 33425 16745 33459 16779
rect 34161 16677 34195 16711
rect 36277 16677 36311 16711
rect 22385 16609 22419 16643
rect 26525 16609 26559 16643
rect 30205 16609 30239 16643
rect 32045 16609 32079 16643
rect 34897 16609 34931 16643
rect 36921 16609 36955 16643
rect 20269 16541 20303 16575
rect 20453 16541 20487 16575
rect 20545 16541 20579 16575
rect 20637 16541 20671 16575
rect 20821 16541 20855 16575
rect 22017 16541 22051 16575
rect 22201 16541 22235 16575
rect 22293 16541 22327 16575
rect 22569 16541 22603 16575
rect 23213 16541 23247 16575
rect 23581 16541 23615 16575
rect 24961 16541 24995 16575
rect 25145 16541 25179 16575
rect 25237 16541 25271 16575
rect 25329 16541 25363 16575
rect 25513 16541 25547 16575
rect 28549 16541 28583 16575
rect 29009 16541 29043 16575
rect 33885 16541 33919 16575
rect 37188 16541 37222 16575
rect 23397 16473 23431 16507
rect 23489 16473 23523 16507
rect 26792 16473 26826 16507
rect 30472 16473 30506 16507
rect 32290 16473 32324 16507
rect 35164 16473 35198 16507
rect 21005 16405 21039 16439
rect 22753 16405 22787 16439
rect 23765 16405 23799 16439
rect 27905 16405 27939 16439
rect 29101 16405 29135 16439
rect 31585 16405 31619 16439
rect 34345 16405 34379 16439
rect 38301 16405 38335 16439
rect 19717 16201 19751 16235
rect 25513 16201 25547 16235
rect 27169 16201 27203 16235
rect 30573 16201 30607 16235
rect 34161 16201 34195 16235
rect 35817 16201 35851 16235
rect 36645 16201 36679 16235
rect 36921 16201 36955 16235
rect 19625 16133 19659 16167
rect 21005 16133 21039 16167
rect 23940 16133 23974 16167
rect 36553 16133 36587 16167
rect 19993 16065 20027 16099
rect 20729 16065 20763 16099
rect 20877 16065 20911 16099
rect 21097 16065 21131 16099
rect 21194 16065 21228 16099
rect 22201 16065 22235 16099
rect 22385 16065 22419 16099
rect 22845 16065 22879 16099
rect 23673 16065 23707 16099
rect 25697 16065 25731 16099
rect 25789 16065 25823 16099
rect 25973 16065 26007 16099
rect 26065 16065 26099 16099
rect 27353 16065 27387 16099
rect 27629 16065 27663 16099
rect 28089 16065 28123 16099
rect 28733 16065 28767 16099
rect 28989 16065 29023 16099
rect 30757 16065 30791 16099
rect 31585 16065 31619 16099
rect 32873 16065 32907 16099
rect 32965 16065 32999 16099
rect 33241 16065 33275 16099
rect 35633 16065 35667 16099
rect 36737 16065 36771 16099
rect 37473 16065 37507 16099
rect 37657 16065 37691 16099
rect 31401 15997 31435 16031
rect 33701 15997 33735 16031
rect 35449 15997 35483 16031
rect 19901 15929 19935 15963
rect 21373 15929 21407 15963
rect 25053 15929 25087 15963
rect 28181 15929 28215 15963
rect 34069 15929 34103 15963
rect 36369 15929 36403 15963
rect 19993 15861 20027 15895
rect 22569 15861 22603 15895
rect 27537 15861 27571 15895
rect 30113 15861 30147 15895
rect 31769 15861 31803 15895
rect 32689 15861 32723 15895
rect 33149 15861 33183 15895
rect 37841 15861 37875 15895
rect 20453 15657 20487 15691
rect 22201 15657 22235 15691
rect 23121 15657 23155 15691
rect 23673 15657 23707 15691
rect 26801 15657 26835 15691
rect 28457 15657 28491 15691
rect 30757 15657 30791 15691
rect 33241 15657 33275 15691
rect 38301 15657 38335 15691
rect 27445 15589 27479 15623
rect 26985 15521 27019 15555
rect 31769 15521 31803 15555
rect 33333 15521 33367 15555
rect 33793 15521 33827 15555
rect 36921 15521 36955 15555
rect 20361 15453 20395 15487
rect 21005 15453 21039 15487
rect 22109 15453 22143 15487
rect 22753 15453 22787 15487
rect 23581 15453 23615 15487
rect 26709 15453 26743 15487
rect 27721 15453 27755 15487
rect 28713 15453 28747 15487
rect 28825 15453 28859 15487
rect 28917 15453 28951 15487
rect 29101 15453 29135 15487
rect 30297 15453 30331 15487
rect 30941 15453 30975 15487
rect 31493 15453 31527 15487
rect 31585 15453 31619 15487
rect 32965 15453 32999 15487
rect 33057 15453 33091 15487
rect 33977 15453 34011 15487
rect 34161 15453 34195 15487
rect 35081 15453 35115 15487
rect 36185 15453 36219 15487
rect 36277 15453 36311 15487
rect 22937 15385 22971 15419
rect 26985 15385 27019 15419
rect 27445 15385 27479 15419
rect 37188 15385 37222 15419
rect 21189 15317 21223 15351
rect 27629 15317 27663 15351
rect 30113 15317 30147 15351
rect 32781 15317 32815 15351
rect 34897 15317 34931 15351
rect 36461 15317 36495 15351
rect 23489 15113 23523 15147
rect 25329 15113 25363 15147
rect 26525 15113 26559 15147
rect 29009 15113 29043 15147
rect 31585 15113 31619 15147
rect 33149 15113 33183 15147
rect 34989 15113 35023 15147
rect 36829 15113 36863 15147
rect 38117 15113 38151 15147
rect 25881 15045 25915 15079
rect 27537 15045 27571 15079
rect 28457 15045 28491 15079
rect 20085 14977 20119 15011
rect 20352 14977 20386 15011
rect 22109 14977 22143 15011
rect 22376 14977 22410 15011
rect 23949 14977 23983 15011
rect 24205 14977 24239 15011
rect 25789 14977 25823 15011
rect 26433 14977 26467 15011
rect 27169 14977 27203 15011
rect 27629 14977 27663 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28917 14977 28951 15011
rect 29101 14977 29135 15011
rect 30461 14977 30495 15011
rect 32965 14977 32999 15011
rect 33609 14977 33643 15011
rect 33876 14977 33910 15011
rect 35449 14977 35483 15011
rect 35705 14977 35739 15011
rect 37657 14977 37691 15011
rect 38301 14977 38335 15011
rect 30205 14909 30239 14943
rect 32781 14909 32815 14943
rect 21465 14773 21499 14807
rect 27353 14773 27387 14807
rect 37473 14773 37507 14807
rect 21281 14569 21315 14603
rect 23397 14569 23431 14603
rect 27629 14569 27663 14603
rect 27813 14569 27847 14603
rect 30021 14569 30055 14603
rect 32597 14569 32631 14603
rect 33057 14569 33091 14603
rect 35265 14569 35299 14603
rect 37289 14569 37323 14603
rect 19441 14433 19475 14467
rect 24961 14433 24995 14467
rect 31217 14433 31251 14467
rect 35909 14433 35943 14467
rect 21557 14365 21591 14399
rect 21646 14362 21680 14396
rect 21741 14359 21775 14393
rect 21925 14365 21959 14399
rect 23673 14365 23707 14399
rect 23762 14359 23796 14393
rect 23862 14365 23896 14399
rect 24041 14365 24075 14399
rect 28457 14365 28491 14399
rect 28641 14365 28675 14399
rect 30205 14365 30239 14399
rect 31473 14365 31507 14399
rect 33057 14365 33091 14399
rect 33241 14365 33275 14399
rect 35449 14365 35483 14399
rect 36176 14365 36210 14399
rect 19708 14297 19742 14331
rect 25228 14297 25262 14331
rect 27445 14297 27479 14331
rect 27661 14297 27695 14331
rect 20821 14229 20855 14263
rect 26341 14229 26375 14263
rect 28641 14229 28675 14263
rect 20453 14025 20487 14059
rect 22937 14025 22971 14059
rect 24041 14025 24075 14059
rect 25145 14025 25179 14059
rect 30205 14025 30239 14059
rect 36185 14025 36219 14059
rect 27721 13957 27755 13991
rect 18889 13889 18923 13923
rect 19717 13889 19751 13923
rect 19901 13889 19935 13923
rect 19993 13889 20027 13923
rect 20085 13889 20119 13923
rect 20280 13889 20314 13923
rect 20913 13889 20947 13923
rect 22201 13889 22235 13923
rect 22385 13889 22419 13923
rect 22569 13889 22603 13923
rect 22753 13889 22787 13923
rect 23765 13889 23799 13923
rect 25421 13889 25455 13923
rect 25513 13889 25547 13923
rect 25605 13889 25639 13923
rect 25789 13889 25823 13923
rect 27905 13889 27939 13923
rect 28825 13889 28859 13923
rect 29092 13889 29126 13923
rect 36001 13889 36035 13923
rect 18981 13821 19015 13855
rect 21189 13821 21223 13855
rect 22477 13821 22511 13855
rect 24041 13821 24075 13855
rect 35817 13821 35851 13855
rect 21005 13753 21039 13787
rect 21097 13753 21131 13787
rect 19165 13685 19199 13719
rect 23857 13685 23891 13719
rect 28089 13685 28123 13719
rect 19993 13481 20027 13515
rect 20545 13481 20579 13515
rect 21281 13481 21315 13515
rect 23029 13481 23063 13515
rect 24961 13481 24995 13515
rect 28549 13481 28583 13515
rect 30113 13481 30147 13515
rect 27997 13413 28031 13447
rect 19625 13345 19659 13379
rect 22385 13345 22419 13379
rect 24685 13345 24719 13379
rect 26249 13345 26283 13379
rect 26985 13345 27019 13379
rect 27721 13345 27755 13379
rect 29745 13345 29779 13379
rect 19809 13277 19843 13311
rect 20453 13277 20487 13311
rect 21189 13277 21223 13311
rect 21373 13277 21407 13311
rect 22753 13277 22787 13311
rect 22845 13277 22879 13311
rect 23489 13277 23523 13311
rect 23673 13277 23707 13311
rect 23949 13277 23983 13311
rect 24961 13277 24995 13311
rect 25145 13277 25179 13311
rect 25973 13277 26007 13311
rect 26065 13277 26099 13311
rect 26709 13277 26743 13311
rect 26801 13277 26835 13311
rect 27629 13277 27663 13311
rect 28779 13277 28813 13311
rect 28917 13277 28951 13311
rect 29030 13277 29064 13311
rect 29193 13277 29227 13311
rect 29929 13277 29963 13311
rect 26985 13209 27019 13243
rect 23857 13141 23891 13175
rect 25605 13141 25639 13175
rect 20085 12937 20119 12971
rect 22385 12937 22419 12971
rect 24133 12937 24167 12971
rect 24685 12937 24719 12971
rect 28273 12937 28307 12971
rect 27353 12869 27387 12903
rect 20269 12801 20303 12835
rect 22293 12801 22327 12835
rect 22477 12801 22511 12835
rect 22937 12801 22971 12835
rect 23029 12801 23063 12835
rect 23949 12801 23983 12835
rect 24593 12801 24627 12835
rect 24777 12801 24811 12835
rect 25421 12801 25455 12835
rect 26249 12801 26283 12835
rect 28181 12801 28215 12835
rect 28365 12801 28399 12835
rect 20545 12733 20579 12767
rect 23213 12733 23247 12767
rect 23765 12733 23799 12767
rect 25329 12733 25363 12767
rect 26525 12733 26559 12767
rect 27629 12733 27663 12767
rect 25789 12665 25823 12699
rect 26341 12665 26375 12699
rect 20453 12597 20487 12631
rect 23121 12597 23155 12631
rect 26433 12597 26467 12631
rect 19809 12393 19843 12427
rect 21373 12393 21407 12427
rect 23029 12393 23063 12427
rect 25973 12393 26007 12427
rect 27353 12393 27387 12427
rect 20913 12325 20947 12359
rect 22569 12325 22603 12359
rect 23305 12325 23339 12359
rect 26341 12325 26375 12359
rect 20637 12257 20671 12291
rect 22109 12257 22143 12291
rect 23397 12257 23431 12291
rect 19717 12189 19751 12223
rect 19901 12189 19935 12223
rect 20545 12189 20579 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 22201 12189 22235 12223
rect 23213 12189 23247 12223
rect 23489 12189 23523 12223
rect 26157 12189 26191 12223
rect 26249 12189 26283 12223
rect 26433 12189 26467 12223
rect 27261 12189 27295 12223
rect 27445 12189 27479 12223
rect 20821 11849 20855 11883
rect 24041 11849 24075 11883
rect 20361 11713 20395 11747
rect 23673 11713 23707 11747
rect 23765 11645 23799 11679
rect 20545 11509 20579 11543
rect 1777 10421 1811 10455
rect 38025 8925 38059 8959
rect 38209 8789 38243 8823
rect 29745 2601 29779 2635
rect 38117 2601 38151 2635
rect 1869 2465 1903 2499
rect 1593 2397 1627 2431
rect 9965 2397 9999 2431
rect 19441 2397 19475 2431
rect 29929 2397 29963 2431
rect 38301 2397 38335 2431
rect 19625 2261 19659 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 29638 37408 29644 37460
rect 29696 37448 29702 37460
rect 29917 37451 29975 37457
rect 29917 37448 29929 37451
rect 29696 37420 29929 37448
rect 29696 37408 29702 37420
rect 29917 37417 29929 37420
rect 29963 37417 29975 37451
rect 29917 37411 29975 37417
rect 38197 37451 38255 37457
rect 38197 37417 38209 37451
rect 38243 37448 38255 37451
rect 39298 37448 39304 37460
rect 38243 37420 39304 37448
rect 38243 37417 38255 37420
rect 38197 37411 38255 37417
rect 39298 37408 39304 37420
rect 39356 37408 39362 37460
rect 658 37204 664 37256
rect 716 37244 722 37256
rect 1765 37247 1823 37253
rect 1765 37244 1777 37247
rect 716 37216 1777 37244
rect 716 37204 722 37216
rect 1765 37213 1777 37216
rect 1811 37213 1823 37247
rect 1765 37207 1823 37213
rect 10318 37204 10324 37256
rect 10376 37244 10382 37256
rect 10505 37247 10563 37253
rect 10505 37244 10517 37247
rect 10376 37216 10517 37244
rect 10376 37204 10382 37216
rect 10505 37213 10517 37216
rect 10551 37213 10563 37247
rect 10505 37207 10563 37213
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20257 37247 20315 37253
rect 20257 37244 20269 37247
rect 20036 37216 20269 37244
rect 20036 37204 20042 37216
rect 20257 37213 20269 37216
rect 20303 37213 20315 37247
rect 20257 37207 20315 37213
rect 32306 37204 32312 37256
rect 32364 37244 32370 37256
rect 38013 37247 38071 37253
rect 38013 37244 38025 37247
rect 32364 37216 38025 37244
rect 32364 37204 32370 37216
rect 38013 37213 38025 37216
rect 38059 37213 38071 37247
rect 38013 37207 38071 37213
rect 1578 37108 1584 37120
rect 1539 37080 1584 37108
rect 1578 37068 1584 37080
rect 1636 37068 1642 37120
rect 10594 37108 10600 37120
rect 10555 37080 10600 37108
rect 10594 37068 10600 37080
rect 10652 37068 10658 37120
rect 20073 37111 20131 37117
rect 20073 37077 20085 37111
rect 20119 37108 20131 37111
rect 24486 37108 24492 37120
rect 20119 37080 24492 37108
rect 20119 37077 20131 37080
rect 20073 37071 20131 37077
rect 24486 37068 24492 37080
rect 24544 37068 24550 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 32306 36904 32312 36916
rect 32267 36876 32312 36904
rect 32306 36864 32312 36876
rect 32364 36864 32370 36916
rect 32490 36768 32496 36780
rect 32451 36740 32496 36768
rect 32490 36728 32496 36740
rect 32548 36728 32554 36780
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 26605 34119 26663 34125
rect 26605 34085 26617 34119
rect 26651 34116 26663 34119
rect 26970 34116 26976 34128
rect 26651 34088 26976 34116
rect 26651 34085 26663 34088
rect 26605 34079 26663 34085
rect 26970 34076 26976 34088
rect 27028 34116 27034 34128
rect 27801 34119 27859 34125
rect 27801 34116 27813 34119
rect 27028 34088 27813 34116
rect 27028 34076 27034 34088
rect 27801 34085 27813 34088
rect 27847 34085 27859 34119
rect 27801 34079 27859 34085
rect 30285 34119 30343 34125
rect 30285 34085 30297 34119
rect 30331 34116 30343 34119
rect 31202 34116 31208 34128
rect 30331 34088 31208 34116
rect 30331 34085 30343 34088
rect 30285 34079 30343 34085
rect 31202 34076 31208 34088
rect 31260 34076 31266 34128
rect 26786 34048 26792 34060
rect 26747 34020 26792 34048
rect 26786 34008 26792 34020
rect 26844 34008 26850 34060
rect 27893 34051 27951 34057
rect 27893 34017 27905 34051
rect 27939 34048 27951 34051
rect 28445 34051 28503 34057
rect 28445 34048 28457 34051
rect 27939 34020 28457 34048
rect 27939 34017 27951 34020
rect 27893 34011 27951 34017
rect 28445 34017 28457 34020
rect 28491 34048 28503 34051
rect 28491 34020 29040 34048
rect 28491 34017 28503 34020
rect 28445 34011 28503 34017
rect 24581 33983 24639 33989
rect 24581 33949 24593 33983
rect 24627 33949 24639 33983
rect 24581 33943 24639 33949
rect 24765 33983 24823 33989
rect 24765 33949 24777 33983
rect 24811 33980 24823 33983
rect 25130 33980 25136 33992
rect 24811 33952 25136 33980
rect 24811 33949 24823 33952
rect 24765 33943 24823 33949
rect 24596 33912 24624 33943
rect 25130 33940 25136 33952
rect 25188 33940 25194 33992
rect 26510 33980 26516 33992
rect 26471 33952 26516 33980
rect 26510 33940 26516 33952
rect 26568 33940 26574 33992
rect 27614 33980 27620 33992
rect 27575 33952 27620 33980
rect 27614 33940 27620 33952
rect 27672 33940 27678 33992
rect 27709 33983 27767 33989
rect 27709 33949 27721 33983
rect 27755 33949 27767 33983
rect 27709 33943 27767 33949
rect 24854 33912 24860 33924
rect 24596 33884 24860 33912
rect 24854 33872 24860 33884
rect 24912 33872 24918 33924
rect 27724 33912 27752 33943
rect 28258 33940 28264 33992
rect 28316 33980 28322 33992
rect 28353 33983 28411 33989
rect 28353 33980 28365 33983
rect 28316 33952 28365 33980
rect 28316 33940 28322 33952
rect 28353 33949 28365 33952
rect 28399 33949 28411 33983
rect 28534 33980 28540 33992
rect 28495 33952 28540 33980
rect 28353 33943 28411 33949
rect 28534 33940 28540 33952
rect 28592 33940 28598 33992
rect 29012 33989 29040 34020
rect 28997 33983 29055 33989
rect 28997 33949 29009 33983
rect 29043 33949 29055 33983
rect 29178 33980 29184 33992
rect 29139 33952 29184 33980
rect 28997 33943 29055 33949
rect 29178 33940 29184 33952
rect 29236 33940 29242 33992
rect 30098 33940 30104 33992
rect 30156 33980 30162 33992
rect 30561 33983 30619 33989
rect 30561 33980 30573 33983
rect 30156 33952 30573 33980
rect 30156 33940 30162 33952
rect 30561 33949 30573 33952
rect 30607 33949 30619 33983
rect 31018 33980 31024 33992
rect 30979 33952 31024 33980
rect 30561 33943 30619 33949
rect 27724 33884 28488 33912
rect 28460 33856 28488 33884
rect 30190 33872 30196 33924
rect 30248 33912 30254 33924
rect 30285 33915 30343 33921
rect 30285 33912 30297 33915
rect 30248 33884 30297 33912
rect 30248 33872 30254 33884
rect 30285 33881 30297 33884
rect 30331 33881 30343 33915
rect 30576 33912 30604 33943
rect 31018 33940 31024 33952
rect 31076 33940 31082 33992
rect 31205 33983 31263 33989
rect 31205 33949 31217 33983
rect 31251 33980 31263 33983
rect 31662 33980 31668 33992
rect 31251 33952 31668 33980
rect 31251 33949 31263 33952
rect 31205 33943 31263 33949
rect 31662 33940 31668 33952
rect 31720 33940 31726 33992
rect 31113 33915 31171 33921
rect 31113 33912 31125 33915
rect 30576 33884 31125 33912
rect 30285 33875 30343 33881
rect 31113 33881 31125 33884
rect 31159 33881 31171 33915
rect 31113 33875 31171 33881
rect 23842 33804 23848 33856
rect 23900 33844 23906 33856
rect 24673 33847 24731 33853
rect 24673 33844 24685 33847
rect 23900 33816 24685 33844
rect 23900 33804 23906 33816
rect 24673 33813 24685 33816
rect 24719 33813 24731 33847
rect 24673 33807 24731 33813
rect 26789 33847 26847 33853
rect 26789 33813 26801 33847
rect 26835 33844 26847 33847
rect 28350 33844 28356 33856
rect 26835 33816 28356 33844
rect 26835 33813 26847 33816
rect 26789 33807 26847 33813
rect 28350 33804 28356 33816
rect 28408 33804 28414 33856
rect 28442 33804 28448 33856
rect 28500 33844 28506 33856
rect 29089 33847 29147 33853
rect 29089 33844 29101 33847
rect 28500 33816 29101 33844
rect 28500 33804 28506 33816
rect 29089 33813 29101 33816
rect 29135 33813 29147 33847
rect 29089 33807 29147 33813
rect 30469 33847 30527 33853
rect 30469 33813 30481 33847
rect 30515 33844 30527 33847
rect 30558 33844 30564 33856
rect 30515 33816 30564 33844
rect 30515 33813 30527 33816
rect 30469 33807 30527 33813
rect 30558 33804 30564 33816
rect 30616 33804 30622 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 24213 33643 24271 33649
rect 24213 33609 24225 33643
rect 24259 33640 24271 33643
rect 26510 33640 26516 33652
rect 24259 33612 24900 33640
rect 26471 33612 26516 33640
rect 24259 33609 24271 33612
rect 24213 33603 24271 33609
rect 24872 33516 24900 33612
rect 26510 33600 26516 33612
rect 26568 33600 26574 33652
rect 27614 33600 27620 33652
rect 27672 33600 27678 33652
rect 30098 33600 30104 33652
rect 30156 33640 30162 33652
rect 31221 33643 31279 33649
rect 31221 33640 31233 33643
rect 30156 33612 31233 33640
rect 30156 33600 30162 33612
rect 31221 33609 31233 33612
rect 31267 33609 31279 33643
rect 31221 33603 31279 33609
rect 27632 33572 27660 33600
rect 29273 33575 29331 33581
rect 27356 33544 28396 33572
rect 23845 33507 23903 33513
rect 23845 33473 23857 33507
rect 23891 33504 23903 33507
rect 24026 33504 24032 33516
rect 23891 33476 24032 33504
rect 23891 33473 23903 33476
rect 23845 33467 23903 33473
rect 24026 33464 24032 33476
rect 24084 33464 24090 33516
rect 24854 33504 24860 33516
rect 24815 33476 24860 33504
rect 24854 33464 24860 33476
rect 24912 33464 24918 33516
rect 26145 33507 26203 33513
rect 26145 33473 26157 33507
rect 26191 33504 26203 33507
rect 27246 33504 27252 33516
rect 26191 33476 27252 33504
rect 26191 33473 26203 33476
rect 26145 33467 26203 33473
rect 27246 33464 27252 33476
rect 27304 33464 27310 33516
rect 27356 33513 27384 33544
rect 27341 33507 27399 33513
rect 27341 33473 27353 33507
rect 27387 33473 27399 33507
rect 27614 33504 27620 33516
rect 27575 33476 27620 33504
rect 27341 33467 27399 33473
rect 27614 33464 27620 33476
rect 27672 33464 27678 33516
rect 28368 33513 28396 33544
rect 29273 33541 29285 33575
rect 29319 33572 29331 33575
rect 30374 33572 30380 33584
rect 29319 33544 30380 33572
rect 29319 33541 29331 33544
rect 29273 33535 29331 33541
rect 30374 33532 30380 33544
rect 30432 33532 30438 33584
rect 31021 33575 31079 33581
rect 31021 33572 31033 33575
rect 30484 33544 31033 33572
rect 28353 33507 28411 33513
rect 28353 33473 28365 33507
rect 28399 33504 28411 33507
rect 30098 33504 30104 33516
rect 28399 33476 28580 33504
rect 30059 33476 30104 33504
rect 28399 33473 28411 33476
rect 28353 33467 28411 33473
rect 23934 33436 23940 33448
rect 23895 33408 23940 33436
rect 23934 33396 23940 33408
rect 23992 33396 23998 33448
rect 24673 33439 24731 33445
rect 24673 33405 24685 33439
rect 24719 33436 24731 33439
rect 26050 33436 26056 33448
rect 24719 33408 25176 33436
rect 26011 33408 26056 33436
rect 24719 33405 24731 33408
rect 24673 33399 24731 33405
rect 25148 33380 25176 33408
rect 26050 33396 26056 33408
rect 26108 33396 26114 33448
rect 27433 33439 27491 33445
rect 27433 33405 27445 33439
rect 27479 33436 27491 33439
rect 28442 33436 28448 33448
rect 27479 33408 28448 33436
rect 27479 33405 27491 33408
rect 27433 33399 27491 33405
rect 28442 33396 28448 33408
rect 28500 33396 28506 33448
rect 28552 33436 28580 33476
rect 30098 33464 30104 33476
rect 30156 33464 30162 33516
rect 30190 33464 30196 33516
rect 30248 33504 30254 33516
rect 30484 33513 30512 33544
rect 31021 33541 31033 33544
rect 31067 33541 31079 33575
rect 31021 33535 31079 33541
rect 30469 33507 30527 33513
rect 30469 33504 30481 33507
rect 30248 33476 30481 33504
rect 30248 33464 30254 33476
rect 30469 33473 30481 33476
rect 30515 33473 30527 33507
rect 30469 33467 30527 33473
rect 30558 33464 30564 33516
rect 30616 33504 30622 33516
rect 30616 33476 30661 33504
rect 30616 33464 30622 33476
rect 30285 33439 30343 33445
rect 30285 33436 30297 33439
rect 28552 33408 30297 33436
rect 30285 33405 30297 33408
rect 30331 33405 30343 33439
rect 30285 33399 30343 33405
rect 33505 33439 33563 33445
rect 33505 33405 33517 33439
rect 33551 33436 33563 33439
rect 34514 33436 34520 33448
rect 33551 33408 34520 33436
rect 33551 33405 33563 33408
rect 33505 33399 33563 33405
rect 34514 33396 34520 33408
rect 34572 33396 34578 33448
rect 23474 33328 23480 33380
rect 23532 33368 23538 33380
rect 25041 33371 25099 33377
rect 25041 33368 25053 33371
rect 23532 33340 25053 33368
rect 23532 33328 23538 33340
rect 25041 33337 25053 33340
rect 25087 33337 25099 33371
rect 25041 33331 25099 33337
rect 25130 33328 25136 33380
rect 25188 33368 25194 33380
rect 27157 33371 27215 33377
rect 27157 33368 27169 33371
rect 25188 33340 27169 33368
rect 25188 33328 25194 33340
rect 27157 33337 27169 33340
rect 27203 33337 27215 33371
rect 27157 33331 27215 33337
rect 27525 33371 27583 33377
rect 27525 33337 27537 33371
rect 27571 33337 27583 33371
rect 27525 33331 27583 33337
rect 28721 33371 28779 33377
rect 28721 33337 28733 33371
rect 28767 33368 28779 33371
rect 29086 33368 29092 33380
rect 28767 33340 29092 33368
rect 28767 33337 28779 33340
rect 28721 33331 28779 33337
rect 26510 33260 26516 33312
rect 26568 33300 26574 33312
rect 27540 33300 27568 33331
rect 29086 33328 29092 33340
rect 29144 33328 29150 33380
rect 33873 33371 33931 33377
rect 33873 33337 33885 33371
rect 33919 33368 33931 33371
rect 34146 33368 34152 33380
rect 33919 33340 34152 33368
rect 33919 33337 33931 33340
rect 33873 33331 33931 33337
rect 34146 33328 34152 33340
rect 34204 33328 34210 33380
rect 26568 33272 27568 33300
rect 26568 33260 26574 33272
rect 28902 33260 28908 33312
rect 28960 33300 28966 33312
rect 29365 33303 29423 33309
rect 29365 33300 29377 33303
rect 28960 33272 29377 33300
rect 28960 33260 28966 33272
rect 29365 33269 29377 33272
rect 29411 33269 29423 33303
rect 29365 33263 29423 33269
rect 30558 33260 30564 33312
rect 30616 33300 30622 33312
rect 31205 33303 31263 33309
rect 31205 33300 31217 33303
rect 30616 33272 31217 33300
rect 30616 33260 30622 33272
rect 31205 33269 31217 33272
rect 31251 33269 31263 33303
rect 31386 33300 31392 33312
rect 31347 33272 31392 33300
rect 31205 33263 31263 33269
rect 31386 33260 31392 33272
rect 31444 33260 31450 33312
rect 33962 33300 33968 33312
rect 33923 33272 33968 33300
rect 33962 33260 33968 33272
rect 34020 33260 34026 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 26697 33099 26755 33105
rect 26697 33065 26709 33099
rect 26743 33096 26755 33099
rect 26786 33096 26792 33108
rect 26743 33068 26792 33096
rect 26743 33065 26755 33068
rect 26697 33059 26755 33065
rect 26786 33056 26792 33068
rect 26844 33056 26850 33108
rect 27614 33056 27620 33108
rect 27672 33096 27678 33108
rect 27709 33099 27767 33105
rect 27709 33096 27721 33099
rect 27672 33068 27721 33096
rect 27672 33056 27678 33068
rect 27709 33065 27721 33068
rect 27755 33065 27767 33099
rect 29178 33096 29184 33108
rect 29139 33068 29184 33096
rect 27709 33059 27767 33065
rect 29178 33056 29184 33068
rect 29236 33056 29242 33108
rect 30558 33056 30564 33108
rect 30616 33096 30622 33108
rect 30745 33099 30803 33105
rect 30745 33096 30757 33099
rect 30616 33068 30757 33096
rect 30616 33056 30622 33068
rect 30745 33065 30757 33068
rect 30791 33065 30803 33099
rect 30745 33059 30803 33065
rect 31297 33099 31355 33105
rect 31297 33065 31309 33099
rect 31343 33096 31355 33099
rect 31386 33096 31392 33108
rect 31343 33068 31392 33096
rect 31343 33065 31355 33068
rect 31297 33059 31355 33065
rect 31386 33056 31392 33068
rect 31444 33056 31450 33108
rect 33962 33096 33968 33108
rect 33923 33068 33968 33096
rect 33962 33056 33968 33068
rect 34020 33056 34026 33108
rect 23474 33028 23480 33040
rect 23032 33000 23480 33028
rect 23032 32901 23060 33000
rect 23474 32988 23480 33000
rect 23532 32988 23538 33040
rect 23750 33028 23756 33040
rect 23711 33000 23756 33028
rect 23750 32988 23756 33000
rect 23808 32988 23814 33040
rect 24854 32988 24860 33040
rect 24912 33028 24918 33040
rect 25225 33031 25283 33037
rect 25225 33028 25237 33031
rect 24912 33000 25237 33028
rect 24912 32988 24918 33000
rect 25225 32997 25237 33000
rect 25271 32997 25283 33031
rect 25225 32991 25283 32997
rect 26528 33000 29776 33028
rect 23293 32963 23351 32969
rect 23293 32929 23305 32963
rect 23339 32960 23351 32963
rect 24578 32960 24584 32972
rect 23339 32932 24584 32960
rect 23339 32929 23351 32932
rect 23293 32923 23351 32929
rect 24578 32920 24584 32932
rect 24636 32960 24642 32972
rect 26528 32969 26556 33000
rect 29748 32972 29776 33000
rect 34514 32988 34520 33040
rect 34572 33028 34578 33040
rect 35161 33031 35219 33037
rect 35161 33028 35173 33031
rect 34572 33000 35173 33028
rect 34572 32988 34578 33000
rect 35161 32997 35173 33000
rect 35207 32997 35219 33031
rect 35161 32991 35219 32997
rect 26513 32963 26571 32969
rect 26513 32960 26525 32963
rect 24636 32932 26525 32960
rect 24636 32920 24642 32932
rect 26513 32929 26525 32932
rect 26559 32929 26571 32963
rect 26513 32923 26571 32929
rect 27801 32963 27859 32969
rect 27801 32929 27813 32963
rect 27847 32960 27859 32963
rect 28258 32960 28264 32972
rect 27847 32932 28264 32960
rect 27847 32929 27859 32932
rect 27801 32923 27859 32929
rect 28258 32920 28264 32932
rect 28316 32960 28322 32972
rect 28902 32960 28908 32972
rect 28316 32932 28908 32960
rect 28316 32920 28322 32932
rect 28902 32920 28908 32932
rect 28960 32920 28966 32972
rect 29730 32920 29736 32972
rect 29788 32960 29794 32972
rect 31481 32963 31539 32969
rect 31481 32960 31493 32963
rect 29788 32932 31493 32960
rect 29788 32920 29794 32932
rect 31481 32929 31493 32932
rect 31527 32960 31539 32963
rect 33505 32963 33563 32969
rect 33505 32960 33517 32963
rect 31527 32932 33517 32960
rect 31527 32929 31539 32932
rect 31481 32923 31539 32929
rect 33505 32929 33517 32932
rect 33551 32929 33563 32963
rect 34054 32960 34060 32972
rect 33967 32932 34060 32960
rect 33505 32923 33563 32929
rect 34054 32920 34060 32932
rect 34112 32960 34118 32972
rect 35345 32963 35403 32969
rect 35345 32960 35357 32963
rect 34112 32932 35357 32960
rect 34112 32920 34118 32932
rect 35345 32929 35357 32932
rect 35391 32929 35403 32963
rect 35345 32923 35403 32929
rect 23017 32895 23075 32901
rect 23017 32861 23029 32895
rect 23063 32861 23075 32895
rect 23017 32855 23075 32861
rect 23109 32895 23167 32901
rect 23109 32861 23121 32895
rect 23155 32892 23167 32895
rect 23753 32895 23811 32901
rect 23753 32892 23765 32895
rect 23155 32864 23765 32892
rect 23155 32861 23167 32864
rect 23109 32855 23167 32861
rect 23753 32861 23765 32864
rect 23799 32892 23811 32895
rect 23842 32892 23848 32904
rect 23799 32864 23848 32892
rect 23799 32861 23811 32864
rect 23753 32855 23811 32861
rect 23842 32852 23848 32864
rect 23900 32852 23906 32904
rect 23934 32852 23940 32904
rect 23992 32892 23998 32904
rect 24029 32895 24087 32901
rect 24029 32892 24041 32895
rect 23992 32864 24041 32892
rect 23992 32852 23998 32864
rect 24029 32861 24041 32864
rect 24075 32892 24087 32895
rect 24854 32892 24860 32904
rect 24075 32864 24860 32892
rect 24075 32861 24087 32864
rect 24029 32855 24087 32861
rect 24854 32852 24860 32864
rect 24912 32852 24918 32904
rect 25130 32892 25136 32904
rect 25091 32864 25136 32892
rect 25130 32852 25136 32864
rect 25188 32852 25194 32904
rect 25222 32852 25228 32904
rect 25280 32892 25286 32904
rect 25317 32895 25375 32901
rect 25317 32892 25329 32895
rect 25280 32864 25329 32892
rect 25280 32852 25286 32864
rect 25317 32861 25329 32864
rect 25363 32861 25375 32895
rect 25317 32855 25375 32861
rect 25409 32895 25467 32901
rect 25409 32861 25421 32895
rect 25455 32892 25467 32895
rect 25958 32892 25964 32904
rect 25455 32864 25964 32892
rect 25455 32861 25467 32864
rect 25409 32855 25467 32861
rect 25958 32852 25964 32864
rect 26016 32852 26022 32904
rect 26970 32892 26976 32904
rect 26931 32864 26976 32892
rect 26970 32852 26976 32864
rect 27028 32852 27034 32904
rect 27246 32852 27252 32904
rect 27304 32892 27310 32904
rect 27525 32895 27583 32901
rect 27525 32892 27537 32895
rect 27304 32864 27537 32892
rect 27304 32852 27310 32864
rect 27525 32861 27537 32864
rect 27571 32861 27583 32895
rect 27525 32855 27583 32861
rect 27617 32895 27675 32901
rect 27617 32861 27629 32895
rect 27663 32861 27675 32895
rect 27617 32855 27675 32861
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 31202 32892 31208 32904
rect 28859 32864 30420 32892
rect 31163 32864 31208 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 23293 32827 23351 32833
rect 23293 32793 23305 32827
rect 23339 32824 23351 32827
rect 25038 32824 25044 32836
rect 23339 32796 25044 32824
rect 23339 32793 23351 32796
rect 23293 32787 23351 32793
rect 25038 32784 25044 32796
rect 25096 32784 25102 32836
rect 27632 32824 27660 32855
rect 30392 32836 30420 32864
rect 31202 32852 31208 32864
rect 31260 32852 31266 32904
rect 33686 32892 33692 32904
rect 33647 32864 33692 32892
rect 33686 32852 33692 32864
rect 33744 32852 33750 32904
rect 33778 32852 33784 32904
rect 33836 32892 33842 32904
rect 33836 32864 33881 32892
rect 33836 32852 33842 32864
rect 28442 32824 28448 32836
rect 27632 32796 28448 32824
rect 28442 32784 28448 32796
rect 28500 32824 28506 32836
rect 28997 32827 29055 32833
rect 28997 32824 29009 32827
rect 28500 32796 29009 32824
rect 28500 32784 28506 32796
rect 28997 32793 29009 32796
rect 29043 32793 29055 32827
rect 30374 32824 30380 32836
rect 30335 32796 30380 32824
rect 28997 32787 29055 32793
rect 30374 32784 30380 32796
rect 30432 32784 30438 32836
rect 30558 32824 30564 32836
rect 30519 32796 30564 32824
rect 30558 32784 30564 32796
rect 30616 32784 30622 32836
rect 34146 32784 34152 32836
rect 34204 32824 34210 32836
rect 34885 32827 34943 32833
rect 34885 32824 34897 32827
rect 34204 32796 34897 32824
rect 34204 32784 34210 32796
rect 34885 32793 34897 32796
rect 34931 32793 34943 32827
rect 34885 32787 34943 32793
rect 23937 32759 23995 32765
rect 23937 32725 23949 32759
rect 23983 32756 23995 32759
rect 24026 32756 24032 32768
rect 23983 32728 24032 32756
rect 23983 32725 23995 32728
rect 23937 32719 23995 32725
rect 24026 32716 24032 32728
rect 24084 32716 24090 32768
rect 24946 32756 24952 32768
rect 24907 32728 24952 32756
rect 24946 32716 24952 32728
rect 25004 32716 25010 32768
rect 26510 32716 26516 32768
rect 26568 32756 26574 32768
rect 26881 32759 26939 32765
rect 26881 32756 26893 32759
rect 26568 32728 26893 32756
rect 26568 32716 26574 32728
rect 26881 32725 26893 32728
rect 26927 32725 26939 32759
rect 26881 32719 26939 32725
rect 30834 32716 30840 32768
rect 30892 32756 30898 32768
rect 31481 32759 31539 32765
rect 31481 32756 31493 32759
rect 30892 32728 31493 32756
rect 30892 32716 30898 32728
rect 31481 32725 31493 32728
rect 31527 32725 31539 32759
rect 31481 32719 31539 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 25222 32552 25228 32564
rect 25183 32524 25228 32552
rect 25222 32512 25228 32524
rect 25280 32512 25286 32564
rect 25958 32552 25964 32564
rect 25919 32524 25964 32552
rect 25958 32512 25964 32524
rect 26016 32512 26022 32564
rect 28442 32552 28448 32564
rect 28276 32524 28448 32552
rect 25240 32484 25268 32512
rect 23860 32456 25268 32484
rect 23860 32425 23888 32456
rect 23845 32419 23903 32425
rect 23845 32385 23857 32419
rect 23891 32385 23903 32419
rect 23845 32379 23903 32385
rect 24857 32419 24915 32425
rect 24857 32385 24869 32419
rect 24903 32416 24915 32419
rect 25130 32416 25136 32428
rect 24903 32388 25136 32416
rect 24903 32385 24915 32388
rect 24857 32379 24915 32385
rect 25130 32376 25136 32388
rect 25188 32416 25194 32428
rect 25685 32419 25743 32425
rect 25685 32416 25697 32419
rect 25188 32388 25697 32416
rect 25188 32376 25194 32388
rect 25685 32385 25697 32388
rect 25731 32385 25743 32419
rect 25685 32379 25743 32385
rect 25774 32376 25780 32428
rect 25832 32416 25838 32428
rect 28166 32416 28172 32428
rect 25832 32388 28172 32416
rect 25832 32376 25838 32388
rect 28166 32376 28172 32388
rect 28224 32376 28230 32428
rect 28276 32425 28304 32524
rect 28442 32512 28448 32524
rect 28500 32512 28506 32564
rect 30374 32512 30380 32564
rect 30432 32552 30438 32564
rect 31018 32552 31024 32564
rect 30432 32524 31024 32552
rect 30432 32512 30438 32524
rect 31018 32512 31024 32524
rect 31076 32552 31082 32564
rect 33413 32555 33471 32561
rect 33413 32552 33425 32555
rect 31076 32524 33425 32552
rect 31076 32512 31082 32524
rect 33413 32521 33425 32524
rect 33459 32521 33471 32555
rect 33778 32552 33784 32564
rect 33413 32515 33471 32521
rect 33612 32524 33784 32552
rect 28368 32456 30696 32484
rect 28368 32425 28396 32456
rect 28261 32419 28319 32425
rect 28261 32385 28273 32419
rect 28307 32385 28319 32419
rect 28261 32379 28319 32385
rect 28353 32419 28411 32425
rect 28353 32385 28365 32419
rect 28399 32385 28411 32419
rect 28353 32379 28411 32385
rect 28445 32419 28503 32425
rect 28445 32385 28457 32419
rect 28491 32385 28503 32419
rect 28626 32416 28632 32428
rect 28587 32388 28632 32416
rect 28445 32379 28503 32385
rect 23750 32348 23756 32360
rect 23711 32320 23756 32348
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 24949 32351 25007 32357
rect 24949 32317 24961 32351
rect 24995 32348 25007 32351
rect 25961 32351 26019 32357
rect 25961 32348 25973 32351
rect 24995 32320 25973 32348
rect 24995 32317 25007 32320
rect 24949 32311 25007 32317
rect 25961 32317 25973 32320
rect 26007 32348 26019 32351
rect 26142 32348 26148 32360
rect 26007 32320 26148 32348
rect 26007 32317 26019 32320
rect 25961 32311 26019 32317
rect 24210 32280 24216 32292
rect 24171 32252 24216 32280
rect 24210 32240 24216 32252
rect 24268 32240 24274 32292
rect 24854 32240 24860 32292
rect 24912 32280 24918 32292
rect 24964 32280 24992 32311
rect 26142 32308 26148 32320
rect 26200 32308 26206 32360
rect 27614 32308 27620 32360
rect 27672 32348 27678 32360
rect 28368 32348 28396 32379
rect 27672 32320 28396 32348
rect 28460 32348 28488 32379
rect 28626 32376 28632 32388
rect 28684 32376 28690 32428
rect 29086 32416 29092 32428
rect 29047 32388 29092 32416
rect 29086 32376 29092 32388
rect 29144 32376 29150 32428
rect 29288 32425 29316 32456
rect 29273 32419 29331 32425
rect 29273 32385 29285 32419
rect 29319 32385 29331 32419
rect 30558 32416 30564 32428
rect 29273 32379 29331 32385
rect 30116 32388 30564 32416
rect 29181 32351 29239 32357
rect 29181 32348 29193 32351
rect 28460 32320 29193 32348
rect 27672 32308 27678 32320
rect 29181 32317 29193 32320
rect 29227 32317 29239 32351
rect 29181 32311 29239 32317
rect 24912 32252 24992 32280
rect 24912 32240 24918 32252
rect 25222 32240 25228 32292
rect 25280 32280 25286 32292
rect 25280 32252 28212 32280
rect 25280 32240 25286 32252
rect 21266 32172 21272 32224
rect 21324 32212 21330 32224
rect 24394 32212 24400 32224
rect 21324 32184 24400 32212
rect 21324 32172 21330 32184
rect 24394 32172 24400 32184
rect 24452 32172 24458 32224
rect 24762 32172 24768 32224
rect 24820 32212 24826 32224
rect 25774 32212 25780 32224
rect 24820 32184 25780 32212
rect 24820 32172 24826 32184
rect 25774 32172 25780 32184
rect 25832 32172 25838 32224
rect 27985 32215 28043 32221
rect 27985 32181 27997 32215
rect 28031 32212 28043 32215
rect 28074 32212 28080 32224
rect 28031 32184 28080 32212
rect 28031 32181 28043 32184
rect 27985 32175 28043 32181
rect 28074 32172 28080 32184
rect 28132 32172 28138 32224
rect 28184 32212 28212 32252
rect 28534 32240 28540 32292
rect 28592 32280 28598 32292
rect 30116 32280 30144 32388
rect 30558 32376 30564 32388
rect 30616 32376 30622 32428
rect 30668 32425 30696 32456
rect 30653 32419 30711 32425
rect 30653 32385 30665 32419
rect 30699 32385 30711 32419
rect 30653 32379 30711 32385
rect 30745 32419 30803 32425
rect 30745 32385 30757 32419
rect 30791 32416 30803 32419
rect 30834 32416 30840 32428
rect 30791 32388 30840 32416
rect 30791 32385 30803 32388
rect 30745 32379 30803 32385
rect 30834 32376 30840 32388
rect 30892 32376 30898 32428
rect 30926 32376 30932 32428
rect 30984 32416 30990 32428
rect 33612 32425 33640 32524
rect 33778 32512 33784 32524
rect 33836 32552 33842 32564
rect 35345 32555 35403 32561
rect 35345 32552 35357 32555
rect 33836 32524 35357 32552
rect 33836 32512 33842 32524
rect 35345 32521 35357 32524
rect 35391 32521 35403 32555
rect 35345 32515 35403 32521
rect 34440 32456 35480 32484
rect 33597 32419 33655 32425
rect 30984 32388 31029 32416
rect 30984 32376 30990 32388
rect 33597 32385 33609 32419
rect 33643 32385 33655 32419
rect 33597 32379 33655 32385
rect 33689 32419 33747 32425
rect 33689 32385 33701 32419
rect 33735 32416 33747 32419
rect 33870 32416 33876 32428
rect 33735 32388 33876 32416
rect 33735 32385 33747 32388
rect 33689 32379 33747 32385
rect 33870 32376 33876 32388
rect 33928 32376 33934 32428
rect 33965 32419 34023 32425
rect 33965 32385 33977 32419
rect 34011 32416 34023 32419
rect 34054 32416 34060 32428
rect 34011 32388 34060 32416
rect 34011 32385 34023 32388
rect 33965 32379 34023 32385
rect 34054 32376 34060 32388
rect 34112 32376 34118 32428
rect 30576 32348 30604 32376
rect 34440 32360 34468 32456
rect 35452 32425 35480 32456
rect 34609 32419 34667 32425
rect 34609 32385 34621 32419
rect 34655 32416 34667 32419
rect 35253 32419 35311 32425
rect 35253 32416 35265 32419
rect 34655 32388 35265 32416
rect 34655 32385 34667 32388
rect 34609 32379 34667 32385
rect 35253 32385 35265 32388
rect 35299 32385 35311 32419
rect 35253 32379 35311 32385
rect 35437 32419 35495 32425
rect 35437 32385 35449 32419
rect 35483 32385 35495 32419
rect 37642 32416 37648 32428
rect 37603 32388 37648 32416
rect 35437 32379 35495 32385
rect 31662 32348 31668 32360
rect 30576 32320 31668 32348
rect 31662 32308 31668 32320
rect 31720 32308 31726 32360
rect 34422 32348 34428 32360
rect 34383 32320 34428 32348
rect 34422 32308 34428 32320
rect 34480 32308 34486 32360
rect 35268 32348 35296 32379
rect 37642 32376 37648 32388
rect 37700 32376 37706 32428
rect 36262 32348 36268 32360
rect 35268 32320 36268 32348
rect 36262 32308 36268 32320
rect 36320 32308 36326 32360
rect 30926 32280 30932 32292
rect 28592 32252 30144 32280
rect 30208 32252 30932 32280
rect 28592 32240 28598 32252
rect 28626 32212 28632 32224
rect 28184 32184 28632 32212
rect 28626 32172 28632 32184
rect 28684 32212 28690 32224
rect 30208 32212 30236 32252
rect 30926 32240 30932 32252
rect 30984 32240 30990 32292
rect 33686 32240 33692 32292
rect 33744 32280 33750 32292
rect 33873 32283 33931 32289
rect 33873 32280 33885 32283
rect 33744 32252 33885 32280
rect 33744 32240 33750 32252
rect 33873 32249 33885 32252
rect 33919 32280 33931 32283
rect 34793 32283 34851 32289
rect 34793 32280 34805 32283
rect 33919 32252 34805 32280
rect 33919 32249 33931 32252
rect 33873 32243 33931 32249
rect 34793 32249 34805 32252
rect 34839 32249 34851 32283
rect 34793 32243 34851 32249
rect 28684 32184 30236 32212
rect 30285 32215 30343 32221
rect 28684 32172 28690 32184
rect 30285 32181 30297 32215
rect 30331 32212 30343 32215
rect 30742 32212 30748 32224
rect 30331 32184 30748 32212
rect 30331 32181 30343 32184
rect 30285 32175 30343 32181
rect 30742 32172 30748 32184
rect 30800 32172 30806 32224
rect 37182 32172 37188 32224
rect 37240 32212 37246 32224
rect 37461 32215 37519 32221
rect 37461 32212 37473 32215
rect 37240 32184 37473 32212
rect 37240 32172 37246 32184
rect 37461 32181 37473 32184
rect 37507 32181 37519 32215
rect 37461 32175 37519 32181
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 21637 32011 21695 32017
rect 21637 31977 21649 32011
rect 21683 32008 21695 32011
rect 31662 32008 31668 32020
rect 21683 31980 31668 32008
rect 21683 31977 21695 31980
rect 21637 31971 21695 31977
rect 31662 31968 31668 31980
rect 31720 31968 31726 32020
rect 31754 31968 31760 32020
rect 31812 32008 31818 32020
rect 32033 32011 32091 32017
rect 32033 32008 32045 32011
rect 31812 31980 32045 32008
rect 31812 31968 31818 31980
rect 32033 31977 32045 31980
rect 32079 31977 32091 32011
rect 32033 31971 32091 31977
rect 33873 32011 33931 32017
rect 33873 31977 33885 32011
rect 33919 32008 33931 32011
rect 34422 32008 34428 32020
rect 33919 31980 34428 32008
rect 33919 31977 33931 31980
rect 33873 31971 33931 31977
rect 34422 31968 34428 31980
rect 34480 31968 34486 32020
rect 36262 32008 36268 32020
rect 36223 31980 36268 32008
rect 36262 31968 36268 31980
rect 36320 31968 36326 32020
rect 23477 31943 23535 31949
rect 23477 31909 23489 31943
rect 23523 31940 23535 31943
rect 24026 31940 24032 31952
rect 23523 31912 24032 31940
rect 23523 31909 23535 31912
rect 23477 31903 23535 31909
rect 24026 31900 24032 31912
rect 24084 31940 24090 31952
rect 24762 31940 24768 31952
rect 24084 31912 24768 31940
rect 24084 31900 24090 31912
rect 24762 31900 24768 31912
rect 24820 31940 24826 31952
rect 24820 31912 24900 31940
rect 24820 31900 24826 31912
rect 21266 31872 21272 31884
rect 21227 31844 21272 31872
rect 21266 31832 21272 31844
rect 21324 31832 21330 31884
rect 21358 31832 21364 31884
rect 21416 31872 21422 31884
rect 22097 31875 22155 31881
rect 22097 31872 22109 31875
rect 21416 31844 22109 31872
rect 21416 31832 21422 31844
rect 22097 31841 22109 31844
rect 22143 31841 22155 31875
rect 22097 31835 22155 31841
rect 24581 31875 24639 31881
rect 24581 31841 24593 31875
rect 24627 31841 24639 31875
rect 24581 31835 24639 31841
rect 1578 31764 1584 31816
rect 1636 31804 1642 31816
rect 20901 31807 20959 31813
rect 20901 31804 20913 31807
rect 1636 31776 20913 31804
rect 1636 31764 1642 31776
rect 20901 31773 20913 31776
rect 20947 31804 20959 31807
rect 21453 31807 21511 31813
rect 21453 31804 21465 31807
rect 20947 31776 21220 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 21192 31736 21220 31776
rect 21376 31776 21465 31804
rect 21376 31736 21404 31776
rect 21453 31773 21465 31776
rect 21499 31773 21511 31807
rect 21453 31767 21511 31773
rect 22364 31807 22422 31813
rect 22364 31773 22376 31807
rect 22410 31804 22422 31807
rect 24596 31804 24624 31835
rect 24872 31813 24900 31912
rect 27246 31900 27252 31952
rect 27304 31940 27310 31952
rect 27430 31940 27436 31952
rect 27304 31912 27436 31940
rect 27304 31900 27310 31912
rect 27430 31900 27436 31912
rect 27488 31940 27494 31952
rect 27488 31912 28212 31940
rect 27488 31900 27494 31912
rect 27893 31875 27951 31881
rect 24964 31844 26004 31872
rect 24964 31813 24992 31844
rect 22410 31776 24624 31804
rect 24857 31807 24915 31813
rect 22410 31773 22422 31776
rect 22364 31767 22422 31773
rect 24857 31773 24869 31807
rect 24903 31773 24915 31807
rect 24857 31767 24915 31773
rect 24949 31807 25007 31813
rect 24949 31773 24961 31807
rect 24995 31773 25007 31807
rect 24949 31767 25007 31773
rect 25038 31764 25044 31816
rect 25096 31804 25102 31816
rect 25222 31804 25228 31816
rect 25096 31776 25141 31804
rect 25183 31776 25228 31804
rect 25096 31764 25102 31776
rect 25222 31764 25228 31776
rect 25280 31764 25286 31816
rect 21192 31708 21404 31736
rect 25976 31736 26004 31844
rect 27893 31841 27905 31875
rect 27939 31841 27951 31875
rect 27893 31835 27951 31841
rect 26050 31764 26056 31816
rect 26108 31804 26114 31816
rect 26320 31807 26378 31813
rect 26108 31776 26153 31804
rect 26108 31764 26114 31776
rect 26320 31773 26332 31807
rect 26366 31804 26378 31807
rect 27908 31804 27936 31835
rect 28184 31813 28212 31912
rect 37274 31900 37280 31952
rect 37332 31940 37338 31952
rect 38105 31943 38163 31949
rect 38105 31940 38117 31943
rect 37332 31912 38117 31940
rect 37332 31900 37338 31912
rect 38105 31909 38117 31912
rect 38151 31909 38163 31943
rect 38105 31903 38163 31909
rect 26366 31776 27936 31804
rect 28169 31807 28227 31813
rect 26366 31773 26378 31776
rect 26320 31767 26378 31773
rect 28169 31773 28181 31807
rect 28215 31773 28227 31807
rect 28169 31767 28227 31773
rect 28261 31807 28319 31813
rect 28261 31773 28273 31807
rect 28307 31773 28319 31807
rect 28261 31767 28319 31773
rect 25976 31708 26280 31736
rect 26252 31680 26280 31708
rect 26602 31696 26608 31748
rect 26660 31736 26666 31748
rect 26660 31708 27292 31736
rect 26660 31696 26666 31708
rect 26234 31628 26240 31680
rect 26292 31628 26298 31680
rect 27264 31668 27292 31708
rect 27614 31696 27620 31748
rect 27672 31736 27678 31748
rect 28276 31736 28304 31767
rect 28350 31764 28356 31816
rect 28408 31804 28414 31816
rect 28537 31807 28595 31813
rect 28408 31776 28453 31804
rect 28408 31764 28414 31776
rect 28537 31773 28549 31807
rect 28583 31804 28595 31807
rect 28626 31804 28632 31816
rect 28583 31776 28632 31804
rect 28583 31773 28595 31776
rect 28537 31767 28595 31773
rect 28626 31764 28632 31776
rect 28684 31764 28690 31816
rect 29730 31804 29736 31816
rect 29691 31776 29736 31804
rect 29730 31764 29736 31776
rect 29788 31764 29794 31816
rect 30653 31807 30711 31813
rect 30653 31773 30665 31807
rect 30699 31773 30711 31807
rect 30653 31767 30711 31773
rect 27672 31708 29960 31736
rect 27672 31696 27678 31708
rect 28902 31668 28908 31680
rect 27264 31640 28908 31668
rect 28902 31628 28908 31640
rect 28960 31628 28966 31680
rect 29932 31677 29960 31708
rect 30282 31696 30288 31748
rect 30340 31736 30346 31748
rect 30668 31736 30696 31767
rect 30742 31764 30748 31816
rect 30800 31804 30806 31816
rect 30909 31807 30967 31813
rect 30909 31804 30921 31807
rect 30800 31776 30921 31804
rect 30800 31764 30806 31776
rect 30909 31773 30921 31776
rect 30955 31773 30967 31807
rect 32490 31804 32496 31816
rect 32451 31776 32496 31804
rect 30909 31767 30967 31773
rect 32490 31764 32496 31776
rect 32548 31764 32554 31816
rect 34606 31764 34612 31816
rect 34664 31804 34670 31816
rect 34885 31807 34943 31813
rect 34664 31776 34836 31804
rect 34664 31764 34670 31776
rect 30340 31708 30696 31736
rect 30340 31696 30346 31708
rect 32398 31696 32404 31748
rect 32456 31736 32462 31748
rect 32738 31739 32796 31745
rect 32738 31736 32750 31739
rect 32456 31708 32750 31736
rect 32456 31696 32462 31708
rect 32738 31705 32750 31708
rect 32784 31705 32796 31739
rect 34808 31736 34836 31776
rect 34885 31773 34897 31807
rect 34931 31804 34943 31807
rect 35526 31804 35532 31816
rect 34931 31776 35532 31804
rect 34931 31773 34943 31776
rect 34885 31767 34943 31773
rect 35526 31764 35532 31776
rect 35584 31764 35590 31816
rect 36906 31804 36912 31816
rect 36867 31776 36912 31804
rect 36906 31764 36912 31776
rect 36964 31764 36970 31816
rect 37645 31807 37703 31813
rect 37645 31773 37657 31807
rect 37691 31804 37703 31807
rect 37826 31804 37832 31816
rect 37691 31776 37832 31804
rect 37691 31773 37703 31776
rect 37645 31767 37703 31773
rect 37826 31764 37832 31776
rect 37884 31764 37890 31816
rect 38286 31804 38292 31816
rect 38247 31776 38292 31804
rect 38286 31764 38292 31776
rect 38344 31764 38350 31816
rect 35130 31739 35188 31745
rect 35130 31736 35142 31739
rect 34808 31708 35142 31736
rect 32738 31699 32796 31705
rect 35130 31705 35142 31708
rect 35176 31705 35188 31739
rect 35130 31699 35188 31705
rect 29917 31671 29975 31677
rect 29917 31637 29929 31671
rect 29963 31668 29975 31671
rect 30098 31668 30104 31680
rect 29963 31640 30104 31668
rect 29963 31637 29975 31640
rect 29917 31631 29975 31637
rect 30098 31628 30104 31640
rect 30156 31628 30162 31680
rect 36722 31668 36728 31680
rect 36683 31640 36728 31668
rect 36722 31628 36728 31640
rect 36780 31628 36786 31680
rect 37458 31668 37464 31680
rect 37419 31640 37464 31668
rect 37458 31628 37464 31640
rect 37516 31628 37522 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 26234 31424 26240 31476
rect 26292 31464 26298 31476
rect 27614 31464 27620 31476
rect 26292 31436 27620 31464
rect 26292 31424 26298 31436
rect 27614 31424 27620 31436
rect 27672 31424 27678 31476
rect 30190 31424 30196 31476
rect 30248 31464 30254 31476
rect 31021 31467 31079 31473
rect 31021 31464 31033 31467
rect 30248 31436 31033 31464
rect 30248 31424 30254 31436
rect 31021 31433 31033 31436
rect 31067 31433 31079 31467
rect 32398 31464 32404 31476
rect 32359 31436 32404 31464
rect 31021 31427 31079 31433
rect 32398 31424 32404 31436
rect 32456 31424 32462 31476
rect 37642 31424 37648 31476
rect 37700 31464 37706 31476
rect 37829 31467 37887 31473
rect 37829 31464 37841 31467
rect 37700 31436 37841 31464
rect 37700 31424 37706 31436
rect 37829 31433 37841 31436
rect 37875 31433 37887 31467
rect 37829 31427 37887 31433
rect 28074 31405 28080 31408
rect 28068 31396 28080 31405
rect 28035 31368 28080 31396
rect 28068 31359 28080 31368
rect 28074 31356 28080 31359
rect 28132 31356 28138 31408
rect 30282 31396 30288 31408
rect 29656 31368 30288 31396
rect 19788 31331 19846 31337
rect 19788 31297 19800 31331
rect 19834 31328 19846 31331
rect 20070 31328 20076 31340
rect 19834 31300 20076 31328
rect 19834 31297 19846 31300
rect 19788 31291 19846 31297
rect 20070 31288 20076 31300
rect 20128 31288 20134 31340
rect 22189 31331 22247 31337
rect 22189 31297 22201 31331
rect 22235 31328 22247 31331
rect 22922 31328 22928 31340
rect 22235 31300 22928 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 22922 31288 22928 31300
rect 22980 31288 22986 31340
rect 26050 31288 26056 31340
rect 26108 31328 26114 31340
rect 27154 31328 27160 31340
rect 26108 31300 27160 31328
rect 26108 31288 26114 31300
rect 27154 31288 27160 31300
rect 27212 31328 27218 31340
rect 29656 31337 29684 31368
rect 30282 31356 30288 31368
rect 30340 31356 30346 31408
rect 33413 31399 33471 31405
rect 33413 31396 33425 31399
rect 32600 31368 33425 31396
rect 27801 31331 27859 31337
rect 27801 31328 27813 31331
rect 27212 31300 27813 31328
rect 27212 31288 27218 31300
rect 27801 31297 27813 31300
rect 27847 31297 27859 31331
rect 27801 31291 27859 31297
rect 29641 31331 29699 31337
rect 29641 31297 29653 31331
rect 29687 31297 29699 31331
rect 29641 31291 29699 31297
rect 29730 31288 29736 31340
rect 29788 31328 29794 31340
rect 29897 31331 29955 31337
rect 29897 31328 29909 31331
rect 29788 31300 29909 31328
rect 29788 31288 29794 31300
rect 29897 31297 29909 31300
rect 29943 31297 29955 31331
rect 31662 31328 31668 31340
rect 31623 31300 31668 31328
rect 29897 31291 29955 31297
rect 31662 31288 31668 31300
rect 31720 31288 31726 31340
rect 32600 31337 32628 31368
rect 33413 31365 33425 31368
rect 33459 31365 33471 31399
rect 33413 31359 33471 31365
rect 35796 31399 35854 31405
rect 35796 31365 35808 31399
rect 35842 31396 35854 31399
rect 36722 31396 36728 31408
rect 35842 31368 36728 31396
rect 35842 31365 35854 31368
rect 35796 31359 35854 31365
rect 36722 31356 36728 31368
rect 36780 31356 36786 31408
rect 32585 31331 32643 31337
rect 32585 31297 32597 31331
rect 32631 31297 32643 31331
rect 33226 31328 33232 31340
rect 33187 31300 33232 31328
rect 32585 31291 32643 31297
rect 33226 31288 33232 31300
rect 33284 31288 33290 31340
rect 35526 31328 35532 31340
rect 35487 31300 35532 31328
rect 35526 31288 35532 31300
rect 35584 31288 35590 31340
rect 36170 31288 36176 31340
rect 36228 31328 36234 31340
rect 37645 31331 37703 31337
rect 37645 31328 37657 31331
rect 36228 31300 37657 31328
rect 36228 31288 36234 31300
rect 37645 31297 37657 31300
rect 37691 31297 37703 31331
rect 37645 31291 37703 31297
rect 19426 31220 19432 31272
rect 19484 31260 19490 31272
rect 19521 31263 19579 31269
rect 19521 31260 19533 31263
rect 19484 31232 19533 31260
rect 19484 31220 19490 31232
rect 19521 31229 19533 31232
rect 19567 31229 19579 31263
rect 19521 31223 19579 31229
rect 22465 31263 22523 31269
rect 22465 31229 22477 31263
rect 22511 31260 22523 31263
rect 22830 31260 22836 31272
rect 22511 31232 22836 31260
rect 22511 31229 22523 31232
rect 22465 31223 22523 31229
rect 22830 31220 22836 31232
rect 22888 31220 22894 31272
rect 33045 31263 33103 31269
rect 33045 31229 33057 31263
rect 33091 31260 33103 31263
rect 34422 31260 34428 31272
rect 33091 31232 34428 31260
rect 33091 31229 33103 31232
rect 33045 31223 33103 31229
rect 34422 31220 34428 31232
rect 34480 31220 34486 31272
rect 37461 31263 37519 31269
rect 37461 31229 37473 31263
rect 37507 31229 37519 31263
rect 37461 31223 37519 31229
rect 20254 31084 20260 31136
rect 20312 31124 20318 31136
rect 20901 31127 20959 31133
rect 20901 31124 20913 31127
rect 20312 31096 20913 31124
rect 20312 31084 20318 31096
rect 20901 31093 20913 31096
rect 20947 31093 20959 31127
rect 20901 31087 20959 31093
rect 21726 31084 21732 31136
rect 21784 31124 21790 31136
rect 22005 31127 22063 31133
rect 22005 31124 22017 31127
rect 21784 31096 22017 31124
rect 21784 31084 21790 31096
rect 22005 31093 22017 31096
rect 22051 31093 22063 31127
rect 22370 31124 22376 31136
rect 22331 31096 22376 31124
rect 22005 31087 22063 31093
rect 22370 31084 22376 31096
rect 22428 31084 22434 31136
rect 28442 31084 28448 31136
rect 28500 31124 28506 31136
rect 29181 31127 29239 31133
rect 29181 31124 29193 31127
rect 28500 31096 29193 31124
rect 28500 31084 28506 31096
rect 29181 31093 29193 31096
rect 29227 31093 29239 31127
rect 29181 31087 29239 31093
rect 31294 31084 31300 31136
rect 31352 31124 31358 31136
rect 31481 31127 31539 31133
rect 31481 31124 31493 31127
rect 31352 31096 31493 31124
rect 31352 31084 31358 31096
rect 31481 31093 31493 31096
rect 31527 31093 31539 31127
rect 31481 31087 31539 31093
rect 36909 31127 36967 31133
rect 36909 31093 36921 31127
rect 36955 31124 36967 31127
rect 37366 31124 37372 31136
rect 36955 31096 37372 31124
rect 36955 31093 36967 31096
rect 36909 31087 36967 31093
rect 37366 31084 37372 31096
rect 37424 31124 37430 31136
rect 37476 31124 37504 31223
rect 37424 31096 37504 31124
rect 37424 31084 37430 31096
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 17313 30923 17371 30929
rect 17313 30889 17325 30923
rect 17359 30920 17371 30923
rect 17402 30920 17408 30932
rect 17359 30892 17408 30920
rect 17359 30889 17371 30892
rect 17313 30883 17371 30889
rect 17402 30880 17408 30892
rect 17460 30880 17466 30932
rect 20346 30880 20352 30932
rect 20404 30920 20410 30932
rect 22462 30920 22468 30932
rect 20404 30892 22468 30920
rect 20404 30880 20410 30892
rect 22462 30880 22468 30892
rect 22520 30880 22526 30932
rect 22830 30920 22836 30932
rect 22791 30892 22836 30920
rect 22830 30880 22836 30892
rect 22888 30880 22894 30932
rect 24946 30880 24952 30932
rect 25004 30920 25010 30932
rect 25498 30920 25504 30932
rect 25004 30892 25504 30920
rect 25004 30880 25010 30892
rect 25498 30880 25504 30892
rect 25556 30920 25562 30932
rect 25593 30923 25651 30929
rect 25593 30920 25605 30923
rect 25556 30892 25605 30920
rect 25556 30880 25562 30892
rect 25593 30889 25605 30892
rect 25639 30889 25651 30923
rect 29730 30920 29736 30932
rect 29691 30892 29736 30920
rect 25593 30883 25651 30889
rect 29730 30880 29736 30892
rect 29788 30880 29794 30932
rect 30098 30920 30104 30932
rect 30059 30892 30104 30920
rect 30098 30880 30104 30892
rect 30156 30880 30162 30932
rect 33226 30880 33232 30932
rect 33284 30920 33290 30932
rect 36170 30920 36176 30932
rect 33284 30892 36176 30920
rect 33284 30880 33290 30892
rect 36170 30880 36176 30892
rect 36228 30880 36234 30932
rect 36357 30923 36415 30929
rect 36357 30889 36369 30923
rect 36403 30920 36415 30923
rect 36906 30920 36912 30932
rect 36403 30892 36912 30920
rect 36403 30889 36415 30892
rect 36357 30883 36415 30889
rect 36906 30880 36912 30892
rect 36964 30880 36970 30932
rect 25685 30855 25743 30861
rect 25685 30821 25697 30855
rect 25731 30852 25743 30855
rect 29362 30852 29368 30864
rect 25731 30824 29368 30852
rect 25731 30821 25743 30824
rect 25685 30815 25743 30821
rect 29362 30812 29368 30824
rect 29420 30812 29426 30864
rect 35526 30812 35532 30864
rect 35584 30852 35590 30864
rect 35584 30824 35894 30852
rect 35584 30812 35590 30824
rect 25774 30784 25780 30796
rect 25735 30756 25780 30784
rect 25774 30744 25780 30756
rect 25832 30744 25838 30796
rect 28977 30787 29035 30793
rect 28977 30753 28989 30787
rect 29023 30784 29035 30787
rect 35866 30784 35894 30824
rect 36906 30784 36912 30796
rect 29023 30756 29960 30784
rect 35866 30756 36912 30784
rect 29023 30753 29035 30756
rect 28977 30747 29035 30753
rect 1578 30716 1584 30728
rect 1539 30688 1584 30716
rect 1578 30676 1584 30688
rect 1636 30676 1642 30728
rect 17034 30716 17040 30728
rect 16995 30688 17040 30716
rect 17034 30676 17040 30688
rect 17092 30676 17098 30728
rect 18598 30676 18604 30728
rect 18656 30716 18662 30728
rect 19429 30719 19487 30725
rect 19429 30716 19441 30719
rect 18656 30688 19441 30716
rect 18656 30676 18662 30688
rect 19429 30685 19441 30688
rect 19475 30685 19487 30719
rect 19429 30679 19487 30685
rect 19613 30719 19671 30725
rect 19613 30685 19625 30719
rect 19659 30685 19671 30719
rect 20254 30716 20260 30728
rect 20215 30688 20260 30716
rect 19613 30679 19671 30685
rect 19628 30648 19656 30679
rect 20254 30676 20260 30688
rect 20312 30676 20318 30728
rect 21358 30676 21364 30728
rect 21416 30716 21422 30728
rect 21453 30719 21511 30725
rect 21453 30716 21465 30719
rect 21416 30688 21465 30716
rect 21416 30676 21422 30688
rect 21453 30685 21465 30688
rect 21499 30716 21511 30719
rect 22002 30716 22008 30728
rect 21499 30688 22008 30716
rect 21499 30685 21511 30688
rect 21453 30679 21511 30685
rect 22002 30676 22008 30688
rect 22060 30676 22066 30728
rect 24578 30716 24584 30728
rect 24539 30688 24584 30716
rect 24578 30676 24584 30688
rect 24636 30676 24642 30728
rect 24765 30719 24823 30725
rect 24765 30685 24777 30719
rect 24811 30716 24823 30719
rect 25038 30716 25044 30728
rect 24811 30688 25044 30716
rect 24811 30685 24823 30688
rect 24765 30679 24823 30685
rect 25038 30676 25044 30688
rect 25096 30676 25102 30728
rect 25501 30719 25559 30725
rect 25501 30685 25513 30719
rect 25547 30685 25559 30719
rect 26234 30716 26240 30728
rect 26195 30688 26240 30716
rect 25501 30679 25559 30685
rect 20162 30648 20168 30660
rect 19628 30620 20168 30648
rect 20162 30608 20168 30620
rect 20220 30608 20226 30660
rect 21726 30657 21732 30660
rect 21720 30648 21732 30657
rect 21687 30620 21732 30648
rect 21720 30611 21732 30620
rect 21726 30608 21732 30611
rect 21784 30608 21790 30660
rect 25516 30648 25544 30679
rect 26234 30676 26240 30688
rect 26292 30676 26298 30728
rect 26421 30719 26479 30725
rect 26421 30685 26433 30719
rect 26467 30716 26479 30719
rect 26602 30716 26608 30728
rect 26467 30688 26608 30716
rect 26467 30685 26479 30688
rect 26421 30679 26479 30685
rect 26602 30676 26608 30688
rect 26660 30676 26666 30728
rect 26878 30716 26884 30728
rect 26839 30688 26884 30716
rect 26878 30676 26884 30688
rect 26936 30676 26942 30728
rect 27065 30719 27123 30725
rect 27065 30685 27077 30719
rect 27111 30716 27123 30719
rect 27614 30716 27620 30728
rect 27111 30688 27620 30716
rect 27111 30685 27123 30688
rect 27065 30679 27123 30685
rect 27614 30676 27620 30688
rect 27672 30676 27678 30728
rect 29178 30716 29184 30728
rect 29091 30688 29184 30716
rect 29178 30676 29184 30688
rect 29236 30716 29242 30728
rect 29638 30716 29644 30728
rect 29236 30688 29644 30716
rect 29236 30676 29242 30688
rect 29638 30676 29644 30688
rect 29696 30676 29702 30728
rect 29932 30725 29960 30756
rect 36906 30744 36912 30756
rect 36964 30744 36970 30796
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30685 29975 30719
rect 30190 30716 30196 30728
rect 30103 30688 30196 30716
rect 29917 30679 29975 30685
rect 30190 30676 30196 30688
rect 30248 30676 30254 30728
rect 30282 30676 30288 30728
rect 30340 30716 30346 30728
rect 31021 30719 31079 30725
rect 31021 30716 31033 30719
rect 30340 30688 31033 30716
rect 30340 30676 30346 30688
rect 31021 30685 31033 30688
rect 31067 30716 31079 30719
rect 32490 30716 32496 30728
rect 31067 30688 32496 30716
rect 31067 30685 31079 30688
rect 31021 30679 31079 30685
rect 25866 30648 25872 30660
rect 25516 30620 25872 30648
rect 25866 30608 25872 30620
rect 25924 30648 25930 30660
rect 26329 30651 26387 30657
rect 26329 30648 26341 30651
rect 25924 30620 26341 30648
rect 25924 30608 25930 30620
rect 26329 30617 26341 30620
rect 26375 30617 26387 30651
rect 26329 30611 26387 30617
rect 28718 30608 28724 30660
rect 28776 30648 28782 30660
rect 28905 30651 28963 30657
rect 28905 30648 28917 30651
rect 28776 30620 28917 30648
rect 28776 30608 28782 30620
rect 28905 30617 28917 30620
rect 28951 30648 28963 30651
rect 28994 30648 29000 30660
rect 28951 30620 29000 30648
rect 28951 30617 28963 30620
rect 28905 30611 28963 30617
rect 28994 30608 29000 30620
rect 29052 30608 29058 30660
rect 30208 30648 30236 30676
rect 31404 30660 31432 30688
rect 32490 30676 32496 30688
rect 32548 30716 32554 30728
rect 32861 30719 32919 30725
rect 32861 30716 32873 30719
rect 32548 30688 32873 30716
rect 32548 30676 32554 30688
rect 32861 30685 32873 30688
rect 32907 30685 32919 30719
rect 32861 30679 32919 30685
rect 35529 30719 35587 30725
rect 35529 30685 35541 30719
rect 35575 30716 35587 30719
rect 35710 30716 35716 30728
rect 35575 30688 35716 30716
rect 35575 30685 35587 30688
rect 35529 30679 35587 30685
rect 35710 30676 35716 30688
rect 35768 30676 35774 30728
rect 35989 30719 36047 30725
rect 35989 30685 36001 30719
rect 36035 30685 36047 30719
rect 36170 30716 36176 30728
rect 36131 30688 36176 30716
rect 35989 30679 36047 30685
rect 31294 30657 31300 30660
rect 31288 30648 31300 30657
rect 29104 30620 30236 30648
rect 31255 30620 31300 30648
rect 1762 30580 1768 30592
rect 1723 30552 1768 30580
rect 1762 30540 1768 30552
rect 1820 30540 1826 30592
rect 17218 30540 17224 30592
rect 17276 30580 17282 30592
rect 17497 30583 17555 30589
rect 17497 30580 17509 30583
rect 17276 30552 17509 30580
rect 17276 30540 17282 30552
rect 17497 30549 17509 30552
rect 17543 30549 17555 30583
rect 17497 30543 17555 30549
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 19797 30583 19855 30589
rect 19797 30580 19809 30583
rect 19392 30552 19809 30580
rect 19392 30540 19398 30552
rect 19797 30549 19809 30552
rect 19843 30549 19855 30583
rect 20346 30580 20352 30592
rect 20307 30552 20352 30580
rect 19797 30543 19855 30549
rect 20346 30540 20352 30552
rect 20404 30540 20410 30592
rect 24673 30583 24731 30589
rect 24673 30549 24685 30583
rect 24719 30580 24731 30583
rect 24854 30580 24860 30592
rect 24719 30552 24860 30580
rect 24719 30549 24731 30552
rect 24673 30543 24731 30549
rect 24854 30540 24860 30552
rect 24912 30540 24918 30592
rect 27065 30583 27123 30589
rect 27065 30549 27077 30583
rect 27111 30580 27123 30583
rect 27246 30580 27252 30592
rect 27111 30552 27252 30580
rect 27111 30549 27123 30552
rect 27065 30543 27123 30549
rect 27246 30540 27252 30552
rect 27304 30540 27310 30592
rect 28810 30540 28816 30592
rect 28868 30580 28874 30592
rect 29104 30589 29132 30620
rect 31288 30611 31300 30620
rect 31294 30608 31300 30611
rect 31352 30608 31358 30660
rect 31386 30608 31392 30660
rect 31444 30608 31450 30660
rect 33128 30651 33186 30657
rect 33128 30617 33140 30651
rect 33174 30648 33186 30651
rect 33962 30648 33968 30660
rect 33174 30620 33968 30648
rect 33174 30617 33186 30620
rect 33128 30611 33186 30617
rect 33962 30608 33968 30620
rect 34020 30608 34026 30660
rect 36004 30648 36032 30679
rect 36170 30676 36176 30688
rect 36228 30676 36234 30728
rect 37182 30725 37188 30728
rect 37176 30716 37188 30725
rect 37143 30688 37188 30716
rect 37176 30679 37188 30688
rect 37182 30676 37188 30679
rect 37240 30676 37246 30728
rect 36262 30648 36268 30660
rect 36004 30620 36268 30648
rect 36262 30608 36268 30620
rect 36320 30608 36326 30660
rect 29089 30583 29147 30589
rect 29089 30580 29101 30583
rect 28868 30552 29101 30580
rect 28868 30540 28874 30552
rect 29089 30549 29101 30552
rect 29135 30549 29147 30583
rect 29089 30543 29147 30549
rect 31846 30540 31852 30592
rect 31904 30580 31910 30592
rect 32401 30583 32459 30589
rect 32401 30580 32413 30583
rect 31904 30552 32413 30580
rect 31904 30540 31910 30552
rect 32401 30549 32413 30552
rect 32447 30549 32459 30583
rect 32401 30543 32459 30549
rect 34054 30540 34060 30592
rect 34112 30580 34118 30592
rect 34241 30583 34299 30589
rect 34241 30580 34253 30583
rect 34112 30552 34253 30580
rect 34112 30540 34118 30552
rect 34241 30549 34253 30552
rect 34287 30549 34299 30583
rect 34241 30543 34299 30549
rect 35345 30583 35403 30589
rect 35345 30549 35357 30583
rect 35391 30580 35403 30583
rect 35618 30580 35624 30592
rect 35391 30552 35624 30580
rect 35391 30549 35403 30552
rect 35345 30543 35403 30549
rect 35618 30540 35624 30552
rect 35676 30540 35682 30592
rect 37918 30540 37924 30592
rect 37976 30580 37982 30592
rect 38289 30583 38347 30589
rect 38289 30580 38301 30583
rect 37976 30552 38301 30580
rect 37976 30540 37982 30552
rect 38289 30549 38301 30552
rect 38335 30549 38347 30583
rect 38289 30543 38347 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 19610 30336 19616 30388
rect 19668 30376 19674 30388
rect 20254 30376 20260 30388
rect 19668 30348 20260 30376
rect 19668 30336 19674 30348
rect 20254 30336 20260 30348
rect 20312 30336 20318 30388
rect 28718 30376 28724 30388
rect 26068 30348 28724 30376
rect 19334 30308 19340 30320
rect 18800 30280 19340 30308
rect 16945 30243 17003 30249
rect 16945 30209 16957 30243
rect 16991 30240 17003 30243
rect 17126 30240 17132 30252
rect 16991 30212 17025 30240
rect 17087 30212 17132 30240
rect 16991 30209 17003 30212
rect 16945 30203 17003 30209
rect 16574 30132 16580 30184
rect 16632 30172 16638 30184
rect 16960 30172 16988 30203
rect 17126 30200 17132 30212
rect 17184 30200 17190 30252
rect 17773 30243 17831 30249
rect 17773 30209 17785 30243
rect 17819 30209 17831 30243
rect 17773 30203 17831 30209
rect 17681 30175 17739 30181
rect 17681 30172 17693 30175
rect 16632 30144 17693 30172
rect 16632 30132 16638 30144
rect 17681 30141 17693 30144
rect 17727 30141 17739 30175
rect 17681 30135 17739 30141
rect 17788 30104 17816 30203
rect 18506 30200 18512 30252
rect 18564 30240 18570 30252
rect 18800 30249 18828 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 19518 30268 19524 30320
rect 19576 30308 19582 30320
rect 20042 30311 20100 30317
rect 20042 30308 20054 30311
rect 19576 30280 20054 30308
rect 19576 30268 19582 30280
rect 20042 30277 20054 30280
rect 20088 30277 20100 30311
rect 20042 30271 20100 30277
rect 22002 30268 22008 30320
rect 22060 30308 22066 30320
rect 26068 30308 26096 30348
rect 28718 30336 28724 30348
rect 28776 30336 28782 30388
rect 28997 30379 29055 30385
rect 28997 30345 29009 30379
rect 29043 30376 29055 30379
rect 29178 30376 29184 30388
rect 29043 30348 29184 30376
rect 29043 30345 29055 30348
rect 28997 30339 29055 30345
rect 29178 30336 29184 30348
rect 29236 30336 29242 30388
rect 33962 30376 33968 30388
rect 33923 30348 33968 30376
rect 33962 30336 33968 30348
rect 34020 30336 34026 30388
rect 35526 30336 35532 30388
rect 35584 30336 35590 30388
rect 36725 30379 36783 30385
rect 36725 30345 36737 30379
rect 36771 30345 36783 30379
rect 36725 30339 36783 30345
rect 37829 30379 37887 30385
rect 37829 30345 37841 30379
rect 37875 30376 37887 30379
rect 37918 30376 37924 30388
rect 37875 30348 37924 30376
rect 37875 30345 37887 30348
rect 37829 30339 37887 30345
rect 22060 30280 23612 30308
rect 22060 30268 22066 30280
rect 18601 30243 18659 30249
rect 18601 30240 18613 30243
rect 18564 30212 18613 30240
rect 18564 30200 18570 30212
rect 18601 30209 18613 30212
rect 18647 30209 18659 30243
rect 18601 30203 18659 30209
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 19153 30243 19211 30249
rect 19153 30209 19165 30243
rect 19199 30209 19211 30243
rect 19153 30203 19211 30209
rect 18874 30172 18880 30184
rect 18835 30144 18880 30172
rect 18874 30132 18880 30144
rect 18932 30132 18938 30184
rect 18969 30175 19027 30181
rect 18969 30141 18981 30175
rect 19015 30172 19027 30175
rect 19058 30172 19064 30184
rect 19015 30144 19064 30172
rect 19015 30141 19027 30144
rect 18969 30135 19027 30141
rect 19058 30132 19064 30144
rect 19116 30132 19122 30184
rect 19168 30172 19196 30203
rect 19426 30200 19432 30252
rect 19484 30240 19490 30252
rect 19797 30243 19855 30249
rect 19797 30240 19809 30243
rect 19484 30212 19809 30240
rect 19484 30200 19490 30212
rect 19797 30209 19809 30212
rect 19843 30240 19855 30243
rect 19886 30240 19892 30252
rect 19843 30212 19892 30240
rect 19843 30209 19855 30212
rect 19797 30203 19855 30209
rect 19886 30200 19892 30212
rect 19944 30200 19950 30252
rect 22462 30240 22468 30252
rect 22423 30212 22468 30240
rect 22462 30200 22468 30212
rect 22520 30200 22526 30252
rect 22830 30240 22836 30252
rect 22791 30212 22836 30240
rect 22830 30200 22836 30212
rect 22888 30200 22894 30252
rect 23584 30249 23612 30280
rect 23676 30280 26096 30308
rect 23569 30243 23627 30249
rect 23569 30209 23581 30243
rect 23615 30209 23627 30243
rect 23569 30203 23627 30209
rect 19610 30172 19616 30184
rect 19168 30144 19616 30172
rect 19610 30132 19616 30144
rect 19668 30132 19674 30184
rect 21910 30132 21916 30184
rect 21968 30172 21974 30184
rect 22005 30175 22063 30181
rect 22005 30172 22017 30175
rect 21968 30144 22017 30172
rect 21968 30132 21974 30144
rect 22005 30141 22017 30144
rect 22051 30141 22063 30175
rect 22186 30172 22192 30184
rect 22147 30144 22192 30172
rect 22005 30135 22063 30141
rect 22186 30132 22192 30144
rect 22244 30132 22250 30184
rect 23474 30132 23480 30184
rect 23532 30172 23538 30184
rect 23676 30172 23704 30280
rect 26234 30268 26240 30320
rect 26292 30308 26298 30320
rect 28902 30308 28908 30320
rect 26292 30280 28908 30308
rect 26292 30268 26298 30280
rect 23836 30243 23894 30249
rect 23836 30209 23848 30243
rect 23882 30240 23894 30243
rect 24946 30240 24952 30252
rect 23882 30212 24952 30240
rect 23882 30209 23894 30212
rect 23836 30203 23894 30209
rect 24946 30200 24952 30212
rect 25004 30200 25010 30252
rect 25593 30243 25651 30249
rect 25593 30209 25605 30243
rect 25639 30240 25651 30243
rect 26050 30240 26056 30252
rect 25639 30212 26056 30240
rect 25639 30209 25651 30212
rect 25593 30203 25651 30209
rect 26050 30200 26056 30212
rect 26108 30200 26114 30252
rect 26436 30249 26464 30280
rect 28902 30268 28908 30280
rect 28960 30268 28966 30320
rect 33686 30268 33692 30320
rect 33744 30308 33750 30320
rect 34333 30311 34391 30317
rect 34333 30308 34345 30311
rect 33744 30280 34345 30308
rect 33744 30268 33750 30280
rect 34333 30277 34345 30280
rect 34379 30277 34391 30311
rect 34333 30271 34391 30277
rect 26421 30243 26479 30249
rect 26421 30209 26433 30243
rect 26467 30209 26479 30243
rect 26421 30203 26479 30209
rect 26602 30200 26608 30252
rect 26660 30240 26666 30252
rect 26970 30240 26976 30252
rect 26660 30212 26976 30240
rect 26660 30200 26666 30212
rect 26970 30200 26976 30212
rect 27028 30200 27034 30252
rect 27154 30240 27160 30252
rect 27115 30212 27160 30240
rect 27154 30200 27160 30212
rect 27212 30200 27218 30252
rect 27430 30249 27436 30252
rect 27424 30203 27436 30249
rect 27488 30240 27494 30252
rect 29362 30240 29368 30252
rect 27488 30212 27524 30240
rect 29323 30212 29368 30240
rect 27430 30200 27436 30203
rect 27488 30200 27494 30212
rect 29362 30200 29368 30212
rect 29420 30200 29426 30252
rect 34146 30240 34152 30252
rect 34107 30212 34152 30240
rect 34146 30200 34152 30212
rect 34204 30200 34210 30252
rect 34241 30243 34299 30249
rect 34241 30209 34253 30243
rect 34287 30209 34299 30243
rect 34241 30203 34299 30209
rect 34471 30243 34529 30249
rect 34471 30209 34483 30243
rect 34517 30240 34529 30243
rect 34790 30240 34796 30252
rect 34517 30212 34796 30240
rect 34517 30209 34529 30212
rect 34471 30203 34529 30209
rect 25498 30172 25504 30184
rect 23532 30144 23704 30172
rect 25459 30144 25504 30172
rect 23532 30132 23538 30144
rect 25498 30132 25504 30144
rect 25556 30132 25562 30184
rect 25774 30132 25780 30184
rect 25832 30172 25838 30184
rect 26513 30175 26571 30181
rect 26513 30172 26525 30175
rect 25832 30144 26525 30172
rect 25832 30132 25838 30144
rect 26513 30141 26525 30144
rect 26559 30141 26571 30175
rect 26513 30135 26571 30141
rect 29454 30132 29460 30184
rect 29512 30172 29518 30184
rect 29512 30144 29557 30172
rect 29512 30132 29518 30144
rect 19794 30104 19800 30116
rect 17788 30076 19800 30104
rect 19794 30064 19800 30076
rect 19852 30064 19858 30116
rect 20806 30064 20812 30116
rect 20864 30104 20870 30116
rect 22097 30107 22155 30113
rect 22097 30104 22109 30107
rect 20864 30076 22109 30104
rect 20864 30064 20870 30076
rect 22097 30073 22109 30076
rect 22143 30073 22155 30107
rect 22097 30067 22155 30073
rect 25961 30107 26019 30113
rect 25961 30073 25973 30107
rect 26007 30104 26019 30107
rect 26878 30104 26884 30116
rect 26007 30076 26884 30104
rect 26007 30073 26019 30076
rect 25961 30067 26019 30073
rect 26878 30064 26884 30076
rect 26936 30064 26942 30116
rect 28537 30107 28595 30113
rect 28537 30073 28549 30107
rect 28583 30104 28595 30107
rect 30006 30104 30012 30116
rect 28583 30076 30012 30104
rect 28583 30073 28595 30076
rect 28537 30067 28595 30073
rect 16945 30039 17003 30045
rect 16945 30005 16957 30039
rect 16991 30036 17003 30039
rect 17402 30036 17408 30048
rect 16991 30008 17408 30036
rect 16991 30005 17003 30008
rect 16945 29999 17003 30005
rect 17402 29996 17408 30008
rect 17460 29996 17466 30048
rect 18046 30036 18052 30048
rect 18007 30008 18052 30036
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 19337 30039 19395 30045
rect 19337 30005 19349 30039
rect 19383 30036 19395 30039
rect 20070 30036 20076 30048
rect 19383 30008 20076 30036
rect 19383 30005 19395 30008
rect 19337 29999 19395 30005
rect 20070 29996 20076 30008
rect 20128 29996 20134 30048
rect 21082 29996 21088 30048
rect 21140 30036 21146 30048
rect 21177 30039 21235 30045
rect 21177 30036 21189 30039
rect 21140 30008 21189 30036
rect 21140 29996 21146 30008
rect 21177 30005 21189 30008
rect 21223 30005 21235 30039
rect 21177 29999 21235 30005
rect 24949 30039 25007 30045
rect 24949 30005 24961 30039
rect 24995 30036 25007 30039
rect 25038 30036 25044 30048
rect 24995 30008 25044 30036
rect 24995 30005 25007 30008
rect 24949 29999 25007 30005
rect 25038 29996 25044 30008
rect 25096 29996 25102 30048
rect 26970 29996 26976 30048
rect 27028 30036 27034 30048
rect 28552 30036 28580 30067
rect 30006 30064 30012 30076
rect 30064 30064 30070 30116
rect 27028 30008 28580 30036
rect 27028 29996 27034 30008
rect 28718 29996 28724 30048
rect 28776 30036 28782 30048
rect 29641 30039 29699 30045
rect 29641 30036 29653 30039
rect 28776 30008 29653 30036
rect 28776 29996 28782 30008
rect 29641 30005 29653 30008
rect 29687 30005 29699 30039
rect 34256 30036 34284 30203
rect 34790 30200 34796 30212
rect 34848 30200 34854 30252
rect 35345 30243 35403 30249
rect 35345 30209 35357 30243
rect 35391 30240 35403 30243
rect 35544 30240 35572 30336
rect 35618 30317 35624 30320
rect 35612 30271 35624 30317
rect 35676 30308 35682 30320
rect 35676 30280 35712 30308
rect 35618 30268 35624 30271
rect 35676 30268 35682 30280
rect 36262 30268 36268 30320
rect 36320 30308 36326 30320
rect 36740 30308 36768 30339
rect 37918 30336 37924 30348
rect 37976 30336 37982 30388
rect 37645 30311 37703 30317
rect 37645 30308 37657 30311
rect 36320 30280 37657 30308
rect 36320 30268 36326 30280
rect 37645 30277 37657 30280
rect 37691 30277 37703 30311
rect 37645 30271 37703 30277
rect 35391 30212 35572 30240
rect 35391 30209 35403 30212
rect 35345 30203 35403 30209
rect 37550 30200 37556 30252
rect 37608 30240 37614 30252
rect 37737 30243 37795 30249
rect 37737 30240 37749 30243
rect 37608 30212 37749 30240
rect 37608 30200 37614 30212
rect 37737 30209 37749 30212
rect 37783 30209 37795 30243
rect 37737 30203 37795 30209
rect 34606 30172 34612 30184
rect 34567 30144 34612 30172
rect 34606 30132 34612 30144
rect 34664 30132 34670 30184
rect 38013 30175 38071 30181
rect 38013 30172 38025 30175
rect 36556 30144 38025 30172
rect 36556 30036 36584 30144
rect 38013 30141 38025 30144
rect 38059 30141 38071 30175
rect 38013 30135 38071 30141
rect 37366 30064 37372 30116
rect 37424 30104 37430 30116
rect 37461 30107 37519 30113
rect 37461 30104 37473 30107
rect 37424 30076 37473 30104
rect 37424 30064 37430 30076
rect 37461 30073 37473 30076
rect 37507 30073 37519 30107
rect 37461 30067 37519 30073
rect 34256 30008 36584 30036
rect 29641 29999 29699 30005
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 16485 29835 16543 29841
rect 16485 29801 16497 29835
rect 16531 29832 16543 29835
rect 17034 29832 17040 29844
rect 16531 29804 17040 29832
rect 16531 29801 16543 29804
rect 16485 29795 16543 29801
rect 17034 29792 17040 29804
rect 17092 29792 17098 29844
rect 18785 29835 18843 29841
rect 18785 29801 18797 29835
rect 18831 29832 18843 29835
rect 18874 29832 18880 29844
rect 18831 29804 18880 29832
rect 18831 29801 18843 29804
rect 18785 29795 18843 29801
rect 18874 29792 18880 29804
rect 18932 29792 18938 29844
rect 19429 29835 19487 29841
rect 19429 29801 19441 29835
rect 19475 29832 19487 29835
rect 19518 29832 19524 29844
rect 19475 29804 19524 29832
rect 19475 29801 19487 29804
rect 19429 29795 19487 29801
rect 19518 29792 19524 29804
rect 19576 29792 19582 29844
rect 19794 29792 19800 29844
rect 19852 29832 19858 29844
rect 20346 29832 20352 29844
rect 19852 29804 20352 29832
rect 19852 29792 19858 29804
rect 20346 29792 20352 29804
rect 20404 29792 20410 29844
rect 22186 29792 22192 29844
rect 22244 29832 22250 29844
rect 22465 29835 22523 29841
rect 22465 29832 22477 29835
rect 22244 29804 22477 29832
rect 22244 29792 22250 29804
rect 22465 29801 22477 29804
rect 22511 29801 22523 29835
rect 22922 29832 22928 29844
rect 22883 29804 22928 29832
rect 22465 29795 22523 29801
rect 22922 29792 22928 29804
rect 22980 29792 22986 29844
rect 24854 29832 24860 29844
rect 24815 29804 24860 29832
rect 24854 29792 24860 29804
rect 24912 29792 24918 29844
rect 24946 29792 24952 29844
rect 25004 29832 25010 29844
rect 25866 29832 25872 29844
rect 25004 29804 25049 29832
rect 25827 29804 25872 29832
rect 25004 29792 25010 29804
rect 25866 29792 25872 29804
rect 25924 29792 25930 29844
rect 26050 29832 26056 29844
rect 26011 29804 26056 29832
rect 26050 29792 26056 29804
rect 26108 29792 26114 29844
rect 26697 29835 26755 29841
rect 26697 29801 26709 29835
rect 26743 29832 26755 29835
rect 27430 29832 27436 29844
rect 26743 29804 27436 29832
rect 26743 29801 26755 29804
rect 26697 29795 26755 29801
rect 27430 29792 27436 29804
rect 27488 29792 27494 29844
rect 29454 29792 29460 29844
rect 29512 29832 29518 29844
rect 30193 29835 30251 29841
rect 30193 29832 30205 29835
rect 29512 29804 30205 29832
rect 29512 29792 29518 29804
rect 30193 29801 30205 29804
rect 30239 29801 30251 29835
rect 30193 29795 30251 29801
rect 34146 29792 34152 29844
rect 34204 29832 34210 29844
rect 34333 29835 34391 29841
rect 34333 29832 34345 29835
rect 34204 29804 34345 29832
rect 34204 29792 34210 29804
rect 34333 29801 34345 29804
rect 34379 29801 34391 29835
rect 34333 29795 34391 29801
rect 34790 29792 34796 29844
rect 34848 29832 34854 29844
rect 35253 29835 35311 29841
rect 35253 29832 35265 29835
rect 34848 29804 35265 29832
rect 34848 29792 34854 29804
rect 35253 29801 35265 29804
rect 35299 29801 35311 29835
rect 36262 29832 36268 29844
rect 36223 29804 36268 29832
rect 35253 29795 35311 29801
rect 36262 29792 36268 29804
rect 36320 29792 36326 29844
rect 37550 29832 37556 29844
rect 36924 29804 37556 29832
rect 17144 29736 18000 29764
rect 17144 29708 17172 29736
rect 17126 29696 17132 29708
rect 16592 29668 17132 29696
rect 16393 29631 16451 29637
rect 16393 29597 16405 29631
rect 16439 29628 16451 29631
rect 16482 29628 16488 29640
rect 16439 29600 16488 29628
rect 16439 29597 16451 29600
rect 16393 29591 16451 29597
rect 16482 29588 16488 29600
rect 16540 29588 16546 29640
rect 16592 29637 16620 29668
rect 17126 29656 17132 29668
rect 17184 29656 17190 29708
rect 17310 29696 17316 29708
rect 17271 29668 17316 29696
rect 17310 29656 17316 29668
rect 17368 29656 17374 29708
rect 17972 29696 18000 29736
rect 18046 29724 18052 29776
rect 18104 29764 18110 29776
rect 18693 29767 18751 29773
rect 18693 29764 18705 29767
rect 18104 29736 18705 29764
rect 18104 29724 18110 29736
rect 18693 29733 18705 29736
rect 18739 29764 18751 29767
rect 20162 29764 20168 29776
rect 18739 29736 20168 29764
rect 18739 29733 18751 29736
rect 18693 29727 18751 29733
rect 20162 29724 20168 29736
rect 20220 29724 20226 29776
rect 21450 29724 21456 29776
rect 21508 29764 21514 29776
rect 21910 29764 21916 29776
rect 21508 29736 21916 29764
rect 21508 29724 21514 29736
rect 21910 29724 21916 29736
rect 21968 29764 21974 29776
rect 28626 29764 28632 29776
rect 21968 29736 24992 29764
rect 21968 29724 21974 29736
rect 24964 29708 24992 29736
rect 27356 29736 28632 29764
rect 18782 29696 18788 29708
rect 17972 29668 18788 29696
rect 18782 29656 18788 29668
rect 18840 29656 18846 29708
rect 18877 29699 18935 29705
rect 18877 29665 18889 29699
rect 18923 29665 18935 29699
rect 20806 29696 20812 29708
rect 18877 29659 18935 29665
rect 18984 29668 20812 29696
rect 16577 29631 16635 29637
rect 16577 29597 16589 29631
rect 16623 29597 16635 29631
rect 17218 29628 17224 29640
rect 17179 29600 17224 29628
rect 16577 29591 16635 29597
rect 17218 29588 17224 29600
rect 17276 29588 17282 29640
rect 18598 29628 18604 29640
rect 18559 29600 18604 29628
rect 18598 29588 18604 29600
rect 18656 29588 18662 29640
rect 18690 29588 18696 29640
rect 18748 29628 18754 29640
rect 18892 29628 18920 29659
rect 18748 29600 18920 29628
rect 18748 29588 18754 29600
rect 1578 29520 1584 29572
rect 1636 29560 1642 29572
rect 1636 29532 18828 29560
rect 1636 29520 1642 29532
rect 17589 29495 17647 29501
rect 17589 29461 17601 29495
rect 17635 29492 17647 29495
rect 18690 29492 18696 29504
rect 17635 29464 18696 29492
rect 17635 29461 17647 29464
rect 17589 29455 17647 29461
rect 18690 29452 18696 29464
rect 18748 29452 18754 29504
rect 18800 29492 18828 29532
rect 18984 29492 19012 29668
rect 20806 29656 20812 29668
rect 20864 29656 20870 29708
rect 21177 29699 21235 29705
rect 21177 29665 21189 29699
rect 21223 29696 21235 29699
rect 21818 29696 21824 29708
rect 21223 29668 21824 29696
rect 21223 29665 21235 29668
rect 21177 29659 21235 29665
rect 21818 29656 21824 29668
rect 21876 29696 21882 29708
rect 22005 29699 22063 29705
rect 22005 29696 22017 29699
rect 21876 29668 22017 29696
rect 21876 29656 21882 29668
rect 22005 29665 22017 29668
rect 22051 29665 22063 29699
rect 22005 29659 22063 29665
rect 22097 29699 22155 29705
rect 22097 29665 22109 29699
rect 22143 29696 22155 29699
rect 24946 29696 24952 29708
rect 22143 29668 22876 29696
rect 24859 29668 24952 29696
rect 22143 29665 22155 29668
rect 22097 29659 22155 29665
rect 22848 29640 22876 29668
rect 24946 29656 24952 29668
rect 25004 29656 25010 29708
rect 19058 29588 19064 29640
rect 19116 29628 19122 29640
rect 19705 29631 19763 29637
rect 19705 29628 19717 29631
rect 19116 29600 19717 29628
rect 19116 29588 19122 29600
rect 18800 29464 19012 29492
rect 19260 29492 19288 29600
rect 19705 29597 19717 29600
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29597 19855 29631
rect 19797 29591 19855 29597
rect 19889 29631 19947 29637
rect 19889 29597 19901 29631
rect 19935 29597 19947 29631
rect 20070 29628 20076 29640
rect 20031 29600 20076 29628
rect 19889 29591 19947 29597
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 19812 29560 19840 29591
rect 19392 29532 19840 29560
rect 19904 29560 19932 29591
rect 20070 29588 20076 29600
rect 20128 29588 20134 29640
rect 21082 29628 21088 29640
rect 20272 29600 21088 29628
rect 20162 29560 20168 29572
rect 19904 29532 20168 29560
rect 19392 29520 19398 29532
rect 20162 29520 20168 29532
rect 20220 29520 20226 29572
rect 20272 29492 20300 29600
rect 21082 29588 21088 29600
rect 21140 29588 21146 29640
rect 21729 29631 21787 29637
rect 21729 29597 21741 29631
rect 21775 29597 21787 29631
rect 21729 29591 21787 29597
rect 21913 29631 21971 29637
rect 21913 29597 21925 29631
rect 21959 29628 21971 29631
rect 22281 29631 22339 29637
rect 21959 29600 22094 29628
rect 21959 29597 21971 29600
rect 21913 29591 21971 29597
rect 19260 29464 20300 29492
rect 21744 29492 21772 29591
rect 22066 29572 22094 29600
rect 22281 29597 22293 29631
rect 22327 29628 22339 29631
rect 22462 29628 22468 29640
rect 22327 29600 22468 29628
rect 22327 29597 22339 29600
rect 22281 29591 22339 29597
rect 22462 29588 22468 29600
rect 22520 29588 22526 29640
rect 22830 29588 22836 29640
rect 22888 29628 22894 29640
rect 23109 29631 23167 29637
rect 23109 29628 23121 29631
rect 22888 29600 23121 29628
rect 22888 29588 22894 29600
rect 23109 29597 23121 29600
rect 23155 29597 23167 29631
rect 23109 29591 23167 29597
rect 23198 29588 23204 29640
rect 23256 29628 23262 29640
rect 23256 29600 23301 29628
rect 23256 29588 23262 29600
rect 24210 29588 24216 29640
rect 24268 29628 24274 29640
rect 24581 29631 24639 29637
rect 24581 29628 24593 29631
rect 24268 29600 24593 29628
rect 24268 29588 24274 29600
rect 24581 29597 24593 29600
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 25593 29631 25651 29637
rect 25593 29597 25605 29631
rect 25639 29628 25651 29631
rect 25774 29628 25780 29640
rect 25639 29600 25780 29628
rect 25639 29597 25651 29600
rect 25593 29591 25651 29597
rect 25774 29588 25780 29600
rect 25832 29588 25838 29640
rect 26970 29628 26976 29640
rect 26931 29600 26976 29628
rect 26970 29588 26976 29600
rect 27028 29588 27034 29640
rect 27065 29631 27123 29637
rect 27065 29597 27077 29631
rect 27111 29597 27123 29631
rect 27065 29591 27123 29597
rect 27157 29631 27215 29637
rect 27157 29597 27169 29631
rect 27203 29628 27215 29631
rect 27246 29628 27252 29640
rect 27203 29600 27252 29628
rect 27203 29597 27215 29600
rect 27157 29591 27215 29597
rect 22066 29532 22100 29572
rect 22094 29520 22100 29532
rect 22152 29520 22158 29572
rect 22925 29563 22983 29569
rect 22925 29529 22937 29563
rect 22971 29560 22983 29563
rect 23474 29560 23480 29572
rect 22971 29532 23480 29560
rect 22971 29529 22983 29532
rect 22925 29523 22983 29529
rect 23474 29520 23480 29532
rect 23532 29520 23538 29572
rect 24673 29563 24731 29569
rect 24673 29529 24685 29563
rect 24719 29560 24731 29563
rect 27080 29560 27108 29591
rect 27246 29588 27252 29600
rect 27304 29588 27310 29640
rect 27356 29637 27384 29736
rect 28626 29724 28632 29736
rect 28684 29764 28690 29776
rect 30558 29764 30564 29776
rect 28684 29736 30564 29764
rect 28684 29724 28690 29736
rect 30558 29724 30564 29736
rect 30616 29724 30622 29776
rect 36924 29764 36952 29804
rect 37550 29792 37556 29804
rect 37608 29832 37614 29844
rect 38289 29835 38347 29841
rect 38289 29832 38301 29835
rect 37608 29804 38301 29832
rect 37608 29792 37614 29804
rect 38289 29801 38301 29804
rect 38335 29801 38347 29835
rect 38289 29795 38347 29801
rect 36188 29736 36952 29764
rect 28718 29696 28724 29708
rect 28679 29668 28724 29696
rect 28718 29656 28724 29668
rect 28776 29656 28782 29708
rect 28902 29656 28908 29708
rect 28960 29696 28966 29708
rect 36188 29705 36216 29736
rect 29825 29699 29883 29705
rect 29825 29696 29837 29699
rect 28960 29668 29837 29696
rect 28960 29656 28966 29668
rect 29825 29665 29837 29668
rect 29871 29665 29883 29699
rect 36173 29699 36231 29705
rect 29825 29659 29883 29665
rect 31864 29668 34008 29696
rect 31864 29640 31892 29668
rect 33980 29640 34008 29668
rect 36173 29665 36185 29699
rect 36219 29665 36231 29699
rect 36906 29696 36912 29708
rect 36867 29668 36912 29696
rect 36173 29659 36231 29665
rect 36906 29656 36912 29668
rect 36964 29656 36970 29708
rect 27341 29631 27399 29637
rect 27341 29597 27353 29631
rect 27387 29597 27399 29631
rect 28442 29628 28448 29640
rect 28403 29600 28448 29628
rect 27341 29591 27399 29597
rect 28442 29588 28448 29600
rect 28500 29588 28506 29640
rect 28626 29628 28632 29640
rect 28587 29600 28632 29628
rect 28626 29588 28632 29600
rect 28684 29588 28690 29640
rect 28813 29631 28871 29637
rect 28813 29597 28825 29631
rect 28859 29597 28871 29631
rect 28813 29591 28871 29597
rect 28997 29631 29055 29637
rect 28997 29597 29009 29631
rect 29043 29628 29055 29631
rect 29917 29631 29975 29637
rect 29917 29628 29929 29631
rect 29043 29600 29929 29628
rect 29043 29597 29055 29600
rect 28997 29591 29055 29597
rect 29917 29597 29929 29600
rect 29963 29628 29975 29631
rect 30926 29628 30932 29640
rect 29963 29600 30932 29628
rect 29963 29597 29975 29600
rect 29917 29591 29975 29597
rect 27614 29560 27620 29572
rect 24719 29532 27620 29560
rect 24719 29529 24731 29532
rect 24673 29523 24731 29529
rect 27614 29520 27620 29532
rect 27672 29560 27678 29572
rect 28828 29560 28856 29591
rect 30926 29588 30932 29600
rect 30984 29588 30990 29640
rect 31846 29628 31852 29640
rect 31807 29600 31852 29628
rect 31846 29588 31852 29600
rect 31904 29588 31910 29640
rect 31941 29631 31999 29637
rect 31941 29597 31953 29631
rect 31987 29628 31999 29631
rect 32214 29628 32220 29640
rect 31987 29600 32220 29628
rect 31987 29597 31999 29600
rect 31941 29591 31999 29597
rect 32214 29588 32220 29600
rect 32272 29588 32278 29640
rect 33962 29628 33968 29640
rect 33875 29600 33968 29628
rect 33962 29588 33968 29600
rect 34020 29588 34026 29640
rect 34057 29631 34115 29637
rect 34057 29597 34069 29631
rect 34103 29628 34115 29631
rect 34514 29628 34520 29640
rect 34103 29600 34520 29628
rect 34103 29597 34115 29600
rect 34057 29591 34115 29597
rect 34514 29588 34520 29600
rect 34572 29588 34578 29640
rect 34885 29631 34943 29637
rect 34885 29597 34897 29631
rect 34931 29628 34943 29631
rect 36265 29631 36323 29637
rect 34931 29600 35894 29628
rect 34931 29597 34943 29600
rect 34885 29591 34943 29597
rect 27672 29532 28856 29560
rect 27672 29520 27678 29532
rect 32766 29520 32772 29572
rect 32824 29560 32830 29572
rect 33781 29563 33839 29569
rect 33781 29560 33793 29563
rect 32824 29532 33793 29560
rect 32824 29520 32830 29532
rect 33781 29529 33793 29532
rect 33827 29529 33839 29563
rect 33781 29523 33839 29529
rect 34238 29520 34244 29572
rect 34296 29560 34302 29572
rect 35069 29563 35127 29569
rect 35069 29560 35081 29563
rect 34296 29532 35081 29560
rect 34296 29520 34302 29532
rect 35069 29529 35081 29532
rect 35115 29529 35127 29563
rect 35069 29523 35127 29529
rect 22278 29492 22284 29504
rect 21744 29464 22284 29492
rect 22278 29452 22284 29464
rect 22336 29452 22342 29504
rect 22370 29452 22376 29504
rect 22428 29492 22434 29504
rect 23198 29492 23204 29504
rect 22428 29464 23204 29492
rect 22428 29452 22434 29464
rect 23198 29452 23204 29464
rect 23256 29452 23262 29504
rect 28442 29452 28448 29504
rect 28500 29492 28506 29504
rect 28902 29492 28908 29504
rect 28500 29464 28908 29492
rect 28500 29452 28506 29464
rect 28902 29452 28908 29464
rect 28960 29452 28966 29504
rect 29181 29495 29239 29501
rect 29181 29461 29193 29495
rect 29227 29492 29239 29495
rect 29638 29492 29644 29504
rect 29227 29464 29644 29492
rect 29227 29461 29239 29464
rect 29181 29455 29239 29461
rect 29638 29452 29644 29464
rect 29696 29452 29702 29504
rect 31754 29452 31760 29504
rect 31812 29492 31818 29504
rect 32125 29495 32183 29501
rect 32125 29492 32137 29495
rect 31812 29464 32137 29492
rect 31812 29452 31818 29464
rect 32125 29461 32137 29464
rect 32171 29461 32183 29495
rect 32125 29455 32183 29461
rect 34146 29452 34152 29504
rect 34204 29492 34210 29504
rect 35866 29492 35894 29600
rect 36265 29597 36277 29631
rect 36311 29597 36323 29631
rect 36265 29591 36323 29597
rect 37176 29631 37234 29637
rect 37176 29597 37188 29631
rect 37222 29628 37234 29631
rect 37458 29628 37464 29640
rect 37222 29600 37464 29628
rect 37222 29597 37234 29600
rect 37176 29591 37234 29597
rect 35986 29560 35992 29572
rect 35947 29532 35992 29560
rect 35986 29520 35992 29532
rect 36044 29520 36050 29572
rect 36280 29560 36308 29591
rect 37458 29588 37464 29600
rect 37516 29588 37522 29640
rect 37366 29560 37372 29572
rect 36280 29532 37372 29560
rect 37366 29520 37372 29532
rect 37424 29520 37430 29572
rect 36449 29495 36507 29501
rect 36449 29492 36461 29495
rect 34204 29464 34249 29492
rect 35866 29464 36461 29492
rect 34204 29452 34210 29464
rect 36449 29461 36461 29464
rect 36495 29461 36507 29495
rect 36449 29455 36507 29461
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 16945 29291 17003 29297
rect 16945 29257 16957 29291
rect 16991 29288 17003 29291
rect 18598 29288 18604 29300
rect 16991 29260 18604 29288
rect 16991 29257 17003 29260
rect 16945 29251 17003 29257
rect 18598 29248 18604 29260
rect 18656 29248 18662 29300
rect 18877 29291 18935 29297
rect 18877 29257 18889 29291
rect 18923 29288 18935 29291
rect 20162 29288 20168 29300
rect 18923 29260 20168 29288
rect 18923 29257 18935 29260
rect 18877 29251 18935 29257
rect 20162 29248 20168 29260
rect 20220 29248 20226 29300
rect 23750 29288 23756 29300
rect 22204 29260 23756 29288
rect 18506 29180 18512 29232
rect 18564 29220 18570 29232
rect 19242 29220 19248 29232
rect 18564 29192 19248 29220
rect 18564 29180 18570 29192
rect 19242 29180 19248 29192
rect 19300 29220 19306 29232
rect 20070 29220 20076 29232
rect 19300 29192 20076 29220
rect 19300 29180 19306 29192
rect 20070 29180 20076 29192
rect 20128 29180 20134 29232
rect 17034 29112 17040 29164
rect 17092 29152 17098 29164
rect 17129 29155 17187 29161
rect 17129 29152 17141 29155
rect 17092 29124 17141 29152
rect 17092 29112 17098 29124
rect 17129 29121 17141 29124
rect 17175 29121 17187 29155
rect 17402 29152 17408 29164
rect 17363 29124 17408 29152
rect 17129 29115 17187 29121
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 18690 29152 18696 29164
rect 18651 29124 18696 29152
rect 18690 29112 18696 29124
rect 18748 29112 18754 29164
rect 18877 29155 18935 29161
rect 18877 29121 18889 29155
rect 18923 29152 18935 29155
rect 19334 29152 19340 29164
rect 18923 29124 19340 29152
rect 18923 29121 18935 29124
rect 18877 29115 18935 29121
rect 19334 29112 19340 29124
rect 19392 29112 19398 29164
rect 22204 29161 22232 29260
rect 23750 29248 23756 29260
rect 23808 29248 23814 29300
rect 25038 29248 25044 29300
rect 25096 29288 25102 29300
rect 27614 29288 27620 29300
rect 25096 29260 27620 29288
rect 25096 29248 25102 29260
rect 27614 29248 27620 29260
rect 27672 29248 27678 29300
rect 28626 29248 28632 29300
rect 28684 29288 28690 29300
rect 28905 29291 28963 29297
rect 28905 29288 28917 29291
rect 28684 29260 28917 29288
rect 28684 29248 28690 29260
rect 28905 29257 28917 29260
rect 28951 29257 28963 29291
rect 30926 29288 30932 29300
rect 30887 29260 30932 29288
rect 28905 29251 28963 29257
rect 30926 29248 30932 29260
rect 30984 29248 30990 29300
rect 34238 29288 34244 29300
rect 34199 29260 34244 29288
rect 34238 29248 34244 29260
rect 34296 29248 34302 29300
rect 35621 29291 35679 29297
rect 35621 29257 35633 29291
rect 35667 29288 35679 29291
rect 35710 29288 35716 29300
rect 35667 29260 35716 29288
rect 35667 29257 35679 29260
rect 35621 29251 35679 29257
rect 35710 29248 35716 29260
rect 35768 29248 35774 29300
rect 37826 29288 37832 29300
rect 37787 29260 37832 29288
rect 37826 29248 37832 29260
rect 37884 29248 37890 29300
rect 22281 29223 22339 29229
rect 22281 29189 22293 29223
rect 22327 29220 22339 29223
rect 23078 29223 23136 29229
rect 23078 29220 23090 29223
rect 22327 29192 23090 29220
rect 22327 29189 22339 29192
rect 22281 29183 22339 29189
rect 23078 29189 23090 29192
rect 23124 29189 23136 29223
rect 23078 29183 23136 29189
rect 25869 29223 25927 29229
rect 25869 29189 25881 29223
rect 25915 29220 25927 29223
rect 28534 29220 28540 29232
rect 25915 29192 26556 29220
rect 25915 29189 25927 29192
rect 25869 29183 25927 29189
rect 22189 29155 22247 29161
rect 22189 29121 22201 29155
rect 22235 29121 22247 29155
rect 22370 29152 22376 29164
rect 22331 29124 22376 29152
rect 22189 29115 22247 29121
rect 22370 29112 22376 29124
rect 22428 29112 22434 29164
rect 25685 29155 25743 29161
rect 25685 29121 25697 29155
rect 25731 29152 25743 29155
rect 25774 29152 25780 29164
rect 25731 29124 25780 29152
rect 25731 29121 25743 29124
rect 25685 29115 25743 29121
rect 25774 29112 25780 29124
rect 25832 29112 25838 29164
rect 25961 29155 26019 29161
rect 25961 29121 25973 29155
rect 26007 29121 26019 29155
rect 26418 29152 26424 29164
rect 26379 29124 26424 29152
rect 25961 29115 26019 29121
rect 19978 29044 19984 29096
rect 20036 29084 20042 29096
rect 22002 29084 22008 29096
rect 20036 29056 22008 29084
rect 20036 29044 20042 29056
rect 22002 29044 22008 29056
rect 22060 29084 22066 29096
rect 22833 29087 22891 29093
rect 22833 29084 22845 29087
rect 22060 29056 22845 29084
rect 22060 29044 22066 29056
rect 22833 29053 22845 29056
rect 22879 29053 22891 29087
rect 25976 29084 26004 29115
rect 26418 29112 26424 29124
rect 26476 29112 26482 29164
rect 26528 29161 26556 29192
rect 28092 29192 28540 29220
rect 28092 29161 28120 29192
rect 28534 29180 28540 29192
rect 28592 29180 28598 29232
rect 29454 29220 29460 29232
rect 28828 29192 29460 29220
rect 26513 29155 26571 29161
rect 26513 29121 26525 29155
rect 26559 29152 26571 29155
rect 27985 29155 28043 29161
rect 27985 29152 27997 29155
rect 26559 29124 27997 29152
rect 26559 29121 26571 29124
rect 26513 29115 26571 29121
rect 27985 29121 27997 29124
rect 28031 29121 28043 29155
rect 27985 29115 28043 29121
rect 28077 29155 28135 29161
rect 28077 29121 28089 29155
rect 28123 29121 28135 29155
rect 28077 29115 28135 29121
rect 27062 29084 27068 29096
rect 25976 29056 27068 29084
rect 22833 29047 22891 29053
rect 27062 29044 27068 29056
rect 27120 29044 27126 29096
rect 28000 29084 28028 29115
rect 28258 29112 28264 29164
rect 28316 29152 28322 29164
rect 28828 29161 28856 29192
rect 29454 29180 29460 29192
rect 29512 29180 29518 29232
rect 30282 29220 30288 29232
rect 29564 29192 30288 29220
rect 28353 29155 28411 29161
rect 28353 29152 28365 29155
rect 28316 29124 28365 29152
rect 28316 29112 28322 29124
rect 28353 29121 28365 29124
rect 28399 29152 28411 29155
rect 28813 29155 28871 29161
rect 28399 29124 28580 29152
rect 28399 29121 28411 29124
rect 28353 29115 28411 29121
rect 28552 29096 28580 29124
rect 28813 29121 28825 29155
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 28997 29155 29055 29161
rect 28997 29121 29009 29155
rect 29043 29152 29055 29155
rect 29362 29152 29368 29164
rect 29043 29124 29368 29152
rect 29043 29121 29055 29124
rect 28997 29115 29055 29121
rect 29362 29112 29368 29124
rect 29420 29112 29426 29164
rect 29564 29161 29592 29192
rect 30282 29180 30288 29192
rect 30340 29180 30346 29232
rect 33781 29223 33839 29229
rect 33781 29189 33793 29223
rect 33827 29220 33839 29223
rect 34146 29220 34152 29232
rect 33827 29192 34152 29220
rect 33827 29189 33839 29192
rect 33781 29183 33839 29189
rect 34146 29180 34152 29192
rect 34204 29180 34210 29232
rect 34330 29180 34336 29232
rect 34388 29220 34394 29232
rect 34388 29192 35894 29220
rect 34388 29180 34394 29192
rect 29549 29155 29607 29161
rect 29549 29121 29561 29155
rect 29595 29121 29607 29155
rect 29549 29115 29607 29121
rect 29638 29112 29644 29164
rect 29696 29152 29702 29164
rect 29805 29155 29863 29161
rect 29805 29152 29817 29155
rect 29696 29124 29817 29152
rect 29696 29112 29702 29124
rect 29805 29121 29817 29124
rect 29851 29121 29863 29155
rect 31754 29152 31760 29164
rect 31715 29124 31760 29152
rect 29805 29115 29863 29121
rect 31754 29112 31760 29124
rect 31812 29112 31818 29164
rect 32766 29152 32772 29164
rect 32727 29124 32772 29152
rect 32766 29112 32772 29124
rect 32824 29112 32830 29164
rect 32858 29112 32864 29164
rect 32916 29152 32922 29164
rect 33226 29152 33232 29164
rect 32916 29124 33232 29152
rect 32916 29112 32922 29124
rect 33226 29112 33232 29124
rect 33284 29112 33290 29164
rect 34057 29155 34115 29161
rect 34057 29152 34069 29155
rect 33336 29124 34069 29152
rect 28442 29084 28448 29096
rect 28000 29056 28448 29084
rect 28442 29044 28448 29056
rect 28500 29044 28506 29096
rect 28534 29044 28540 29096
rect 28592 29044 28598 29096
rect 32784 29084 32812 29112
rect 33336 29084 33364 29124
rect 34057 29121 34069 29124
rect 34103 29121 34115 29155
rect 35342 29152 35348 29164
rect 35303 29124 35348 29152
rect 34057 29115 34115 29121
rect 35342 29112 35348 29124
rect 35400 29112 35406 29164
rect 35437 29155 35495 29161
rect 35437 29121 35449 29155
rect 35483 29121 35495 29155
rect 35866 29152 35894 29192
rect 35986 29180 35992 29232
rect 36044 29220 36050 29232
rect 37918 29220 37924 29232
rect 36044 29192 37924 29220
rect 36044 29180 36050 29192
rect 36357 29155 36415 29161
rect 36357 29152 36369 29155
rect 35866 29124 36369 29152
rect 35437 29115 35495 29121
rect 36357 29121 36369 29124
rect 36403 29121 36415 29155
rect 36357 29115 36415 29121
rect 36541 29155 36599 29161
rect 36541 29121 36553 29155
rect 36587 29152 36599 29155
rect 37274 29152 37280 29164
rect 36587 29124 37280 29152
rect 36587 29121 36599 29124
rect 36541 29115 36599 29121
rect 32784 29056 33364 29084
rect 33965 29087 34023 29093
rect 33965 29053 33977 29087
rect 34011 29084 34023 29087
rect 34514 29084 34520 29096
rect 34011 29056 34520 29084
rect 34011 29053 34023 29056
rect 33965 29047 34023 29053
rect 34514 29044 34520 29056
rect 34572 29084 34578 29096
rect 35360 29084 35388 29112
rect 34572 29056 35388 29084
rect 35452 29084 35480 29115
rect 37274 29112 37280 29124
rect 37332 29112 37338 29164
rect 37568 29161 37596 29192
rect 37918 29180 37924 29192
rect 37976 29180 37982 29232
rect 37553 29155 37611 29161
rect 37553 29121 37565 29155
rect 37599 29121 37611 29155
rect 37553 29115 37611 29121
rect 37642 29112 37648 29164
rect 37700 29152 37706 29164
rect 37700 29124 37793 29152
rect 37700 29112 37706 29124
rect 37752 29084 37780 29124
rect 35452 29056 37780 29084
rect 34572 29044 34578 29056
rect 17310 29016 17316 29028
rect 17271 28988 17316 29016
rect 17310 28976 17316 28988
rect 17368 28976 17374 29028
rect 27430 28976 27436 29028
rect 27488 29016 27494 29028
rect 28261 29019 28319 29025
rect 28261 29016 28273 29019
rect 27488 28988 28273 29016
rect 27488 28976 27494 28988
rect 28261 28985 28273 28988
rect 28307 28985 28319 29019
rect 28261 28979 28319 28985
rect 33045 29019 33103 29025
rect 33045 28985 33057 29019
rect 33091 29016 33103 29019
rect 33410 29016 33416 29028
rect 33091 28988 33416 29016
rect 33091 28985 33103 28988
rect 33045 28979 33103 28985
rect 33410 28976 33416 28988
rect 33468 28976 33474 29028
rect 33502 28976 33508 29028
rect 33560 29016 33566 29028
rect 35452 29016 35480 29056
rect 33560 28988 35480 29016
rect 33560 28976 33566 28988
rect 23566 28908 23572 28960
rect 23624 28948 23630 28960
rect 24213 28951 24271 28957
rect 24213 28948 24225 28951
rect 23624 28920 24225 28948
rect 23624 28908 23630 28920
rect 24213 28917 24225 28920
rect 24259 28917 24271 28951
rect 25682 28948 25688 28960
rect 25643 28920 25688 28948
rect 24213 28911 24271 28917
rect 25682 28908 25688 28920
rect 25740 28908 25746 28960
rect 27798 28948 27804 28960
rect 27759 28920 27804 28948
rect 27798 28908 27804 28920
rect 27856 28908 27862 28960
rect 31573 28951 31631 28957
rect 31573 28917 31585 28951
rect 31619 28948 31631 28951
rect 31662 28948 31668 28960
rect 31619 28920 31668 28948
rect 31619 28917 31631 28920
rect 31573 28911 31631 28917
rect 31662 28908 31668 28920
rect 31720 28908 31726 28960
rect 33962 28948 33968 28960
rect 33923 28920 33968 28948
rect 33962 28908 33968 28920
rect 34020 28908 34026 28960
rect 36170 28908 36176 28960
rect 36228 28948 36234 28960
rect 36725 28951 36783 28957
rect 36725 28948 36737 28951
rect 36228 28920 36737 28948
rect 36228 28908 36234 28920
rect 36725 28917 36737 28920
rect 36771 28917 36783 28951
rect 36725 28911 36783 28917
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 22278 28744 22284 28756
rect 22239 28716 22284 28744
rect 22278 28704 22284 28716
rect 22336 28704 22342 28756
rect 22646 28704 22652 28756
rect 22704 28744 22710 28756
rect 22925 28747 22983 28753
rect 22925 28744 22937 28747
rect 22704 28716 22937 28744
rect 22704 28704 22710 28716
rect 22925 28713 22937 28716
rect 22971 28713 22983 28747
rect 22925 28707 22983 28713
rect 23109 28747 23167 28753
rect 23109 28713 23121 28747
rect 23155 28744 23167 28747
rect 23198 28744 23204 28756
rect 23155 28716 23204 28744
rect 23155 28713 23167 28716
rect 23109 28707 23167 28713
rect 23198 28704 23204 28716
rect 23256 28704 23262 28756
rect 23750 28744 23756 28756
rect 23711 28716 23756 28744
rect 23750 28704 23756 28716
rect 23808 28704 23814 28756
rect 24394 28704 24400 28756
rect 24452 28744 24458 28756
rect 26418 28744 26424 28756
rect 24452 28716 26280 28744
rect 26379 28716 26424 28744
rect 24452 28704 24458 28716
rect 22738 28676 22744 28688
rect 21652 28648 22744 28676
rect 19797 28543 19855 28549
rect 19797 28509 19809 28543
rect 19843 28540 19855 28543
rect 19886 28540 19892 28552
rect 19843 28512 19892 28540
rect 19843 28509 19855 28512
rect 19797 28503 19855 28509
rect 19886 28500 19892 28512
rect 19944 28500 19950 28552
rect 21652 28549 21680 28648
rect 22738 28636 22744 28648
rect 22796 28636 22802 28688
rect 26252 28676 26280 28716
rect 26418 28704 26424 28716
rect 26476 28704 26482 28756
rect 30745 28747 30803 28753
rect 30745 28713 30757 28747
rect 30791 28713 30803 28747
rect 30745 28707 30803 28713
rect 30929 28747 30987 28753
rect 30929 28713 30941 28747
rect 30975 28744 30987 28747
rect 32306 28744 32312 28756
rect 30975 28716 32312 28744
rect 30975 28713 30987 28716
rect 30929 28707 30987 28713
rect 29270 28676 29276 28688
rect 26252 28648 29276 28676
rect 29270 28636 29276 28648
rect 29328 28636 29334 28688
rect 30760 28620 30788 28707
rect 32306 28704 32312 28716
rect 32364 28704 32370 28756
rect 32766 28744 32772 28756
rect 32727 28716 32772 28744
rect 32766 28704 32772 28716
rect 32824 28704 32830 28756
rect 35526 28704 35532 28756
rect 35584 28744 35590 28756
rect 38105 28747 38163 28753
rect 38105 28744 38117 28747
rect 35584 28716 38117 28744
rect 35584 28704 35590 28716
rect 38105 28713 38117 28716
rect 38151 28713 38163 28747
rect 38105 28707 38163 28713
rect 21910 28568 21916 28620
rect 21968 28568 21974 28620
rect 23845 28611 23903 28617
rect 22756 28580 23244 28608
rect 21818 28549 21824 28552
rect 21637 28543 21695 28549
rect 21637 28509 21649 28543
rect 21683 28509 21695 28543
rect 21637 28503 21695 28509
rect 21785 28543 21824 28549
rect 21785 28509 21797 28543
rect 21785 28503 21824 28509
rect 21818 28500 21824 28503
rect 21876 28500 21882 28552
rect 21928 28540 21956 28568
rect 22186 28549 22192 28552
rect 22013 28543 22071 28549
rect 22013 28540 22025 28543
rect 21928 28512 22025 28540
rect 22013 28509 22025 28512
rect 22059 28509 22071 28543
rect 22013 28503 22071 28509
rect 22143 28543 22192 28549
rect 22143 28509 22155 28543
rect 22189 28509 22192 28543
rect 22143 28503 22192 28509
rect 22186 28500 22192 28503
rect 22244 28540 22250 28552
rect 22756 28540 22784 28580
rect 22244 28512 22784 28540
rect 22244 28500 22250 28512
rect 20064 28475 20122 28481
rect 20064 28441 20076 28475
rect 20110 28472 20122 28475
rect 20162 28472 20168 28484
rect 20110 28444 20168 28472
rect 20110 28441 20122 28444
rect 20064 28435 20122 28441
rect 20162 28432 20168 28444
rect 20220 28432 20226 28484
rect 21913 28475 21971 28481
rect 21913 28441 21925 28475
rect 21959 28472 21971 28475
rect 22646 28472 22652 28484
rect 21959 28444 22652 28472
rect 21959 28441 21971 28444
rect 21913 28435 21971 28441
rect 22646 28432 22652 28444
rect 22704 28432 22710 28484
rect 22756 28481 22784 28512
rect 23106 28500 23112 28552
rect 23164 28500 23170 28552
rect 23216 28540 23244 28580
rect 23845 28577 23857 28611
rect 23891 28608 23903 28611
rect 24854 28608 24860 28620
rect 23891 28580 24860 28608
rect 23891 28577 23903 28580
rect 23845 28571 23903 28577
rect 24854 28568 24860 28580
rect 24912 28568 24918 28620
rect 30742 28608 30748 28620
rect 28184 28580 30748 28608
rect 23566 28540 23572 28552
rect 23216 28512 23572 28540
rect 23566 28500 23572 28512
rect 23624 28500 23630 28552
rect 23658 28500 23664 28552
rect 23716 28540 23722 28552
rect 25041 28543 25099 28549
rect 23716 28512 23761 28540
rect 23716 28500 23722 28512
rect 25041 28509 25053 28543
rect 25087 28540 25099 28543
rect 26234 28540 26240 28552
rect 25087 28512 26240 28540
rect 25087 28509 25099 28512
rect 25041 28503 25099 28509
rect 26234 28500 26240 28512
rect 26292 28540 26298 28552
rect 27154 28540 27160 28552
rect 26292 28512 27160 28540
rect 26292 28500 26298 28512
rect 27154 28500 27160 28512
rect 27212 28500 27218 28552
rect 27246 28500 27252 28552
rect 27304 28540 27310 28552
rect 27525 28543 27583 28549
rect 27304 28512 27349 28540
rect 27304 28500 27310 28512
rect 27525 28509 27537 28543
rect 27571 28540 27583 28543
rect 28074 28540 28080 28552
rect 27571 28512 28080 28540
rect 27571 28509 27583 28512
rect 27525 28503 27583 28509
rect 28074 28500 28080 28512
rect 28132 28500 28138 28552
rect 28184 28549 28212 28580
rect 30742 28568 30748 28580
rect 30800 28568 30806 28620
rect 33873 28611 33931 28617
rect 33873 28577 33885 28611
rect 33919 28608 33931 28611
rect 34146 28608 34152 28620
rect 33919 28580 34152 28608
rect 33919 28577 33931 28580
rect 33873 28571 33931 28577
rect 34146 28568 34152 28580
rect 34204 28568 34210 28620
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28509 28227 28543
rect 28169 28503 28227 28509
rect 28258 28500 28264 28552
rect 28316 28540 28322 28552
rect 28445 28543 28503 28549
rect 28445 28540 28457 28543
rect 28316 28512 28457 28540
rect 28316 28500 28322 28512
rect 28445 28509 28457 28512
rect 28491 28509 28503 28543
rect 28445 28503 28503 28509
rect 28629 28543 28687 28549
rect 28629 28509 28641 28543
rect 28675 28540 28687 28543
rect 28810 28540 28816 28552
rect 28675 28512 28816 28540
rect 28675 28509 28687 28512
rect 28629 28503 28687 28509
rect 22741 28475 22799 28481
rect 22741 28441 22753 28475
rect 22787 28441 22799 28475
rect 22741 28435 22799 28441
rect 22957 28475 23015 28481
rect 22957 28441 22969 28475
rect 23003 28472 23015 28475
rect 23124 28472 23152 28500
rect 23003 28444 23152 28472
rect 25308 28475 25366 28481
rect 23003 28441 23015 28444
rect 22957 28435 23015 28441
rect 25308 28441 25320 28475
rect 25354 28472 25366 28475
rect 25682 28472 25688 28484
rect 25354 28444 25688 28472
rect 25354 28441 25366 28444
rect 25308 28435 25366 28441
rect 25682 28432 25688 28444
rect 25740 28432 25746 28484
rect 27433 28475 27491 28481
rect 27433 28441 27445 28475
rect 27479 28472 27491 28475
rect 27798 28472 27804 28484
rect 27479 28444 27804 28472
rect 27479 28441 27491 28444
rect 27433 28435 27491 28441
rect 27798 28432 27804 28444
rect 27856 28432 27862 28484
rect 27890 28432 27896 28484
rect 27948 28472 27954 28484
rect 28644 28472 28672 28503
rect 28810 28500 28816 28512
rect 28868 28500 28874 28552
rect 29917 28543 29975 28549
rect 29917 28509 29929 28543
rect 29963 28540 29975 28543
rect 31018 28540 31024 28552
rect 29963 28512 31024 28540
rect 29963 28509 29975 28512
rect 29917 28503 29975 28509
rect 31018 28500 31024 28512
rect 31076 28500 31082 28552
rect 31386 28540 31392 28552
rect 31299 28512 31392 28540
rect 31386 28500 31392 28512
rect 31444 28500 31450 28552
rect 31662 28549 31668 28552
rect 31656 28540 31668 28549
rect 31623 28512 31668 28540
rect 31656 28503 31668 28512
rect 31662 28500 31668 28503
rect 31720 28500 31726 28552
rect 33410 28540 33416 28552
rect 33371 28512 33416 28540
rect 33410 28500 33416 28512
rect 33468 28500 33474 28552
rect 34057 28543 34115 28549
rect 34057 28509 34069 28543
rect 34103 28540 34115 28543
rect 34330 28540 34336 28552
rect 34103 28512 34336 28540
rect 34103 28509 34115 28512
rect 34057 28503 34115 28509
rect 27948 28444 28672 28472
rect 30561 28475 30619 28481
rect 27948 28432 27954 28444
rect 30561 28441 30573 28475
rect 30607 28472 30619 28475
rect 31294 28472 31300 28484
rect 30607 28444 31300 28472
rect 30607 28441 30619 28444
rect 30561 28435 30619 28441
rect 31294 28432 31300 28444
rect 31352 28432 31358 28484
rect 31404 28472 31432 28500
rect 32030 28472 32036 28484
rect 31404 28444 32036 28472
rect 32030 28432 32036 28444
rect 32088 28432 32094 28484
rect 32214 28432 32220 28484
rect 32272 28472 32278 28484
rect 34072 28472 34100 28503
rect 34330 28500 34336 28512
rect 34388 28500 34394 28552
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28540 34943 28543
rect 36725 28543 36783 28549
rect 36725 28540 36737 28543
rect 34931 28512 36737 28540
rect 34931 28509 34943 28512
rect 34885 28503 34943 28509
rect 36725 28509 36737 28512
rect 36771 28540 36783 28543
rect 36814 28540 36820 28552
rect 36771 28512 36820 28540
rect 36771 28509 36783 28512
rect 36725 28503 36783 28509
rect 36814 28500 36820 28512
rect 36872 28500 36878 28552
rect 32272 28444 34100 28472
rect 32272 28432 32278 28444
rect 34790 28432 34796 28484
rect 34848 28472 34854 28484
rect 35130 28475 35188 28481
rect 35130 28472 35142 28475
rect 34848 28444 35142 28472
rect 34848 28432 34854 28444
rect 35130 28441 35142 28444
rect 35176 28441 35188 28475
rect 35130 28435 35188 28441
rect 35986 28432 35992 28484
rect 36044 28472 36050 28484
rect 36970 28475 37028 28481
rect 36970 28472 36982 28475
rect 36044 28444 36982 28472
rect 36044 28432 36050 28444
rect 36970 28441 36982 28444
rect 37016 28441 37028 28475
rect 36970 28435 37028 28441
rect 21174 28404 21180 28416
rect 21135 28376 21180 28404
rect 21174 28364 21180 28376
rect 21232 28364 21238 28416
rect 21818 28364 21824 28416
rect 21876 28404 21882 28416
rect 22094 28404 22100 28416
rect 21876 28376 22100 28404
rect 21876 28364 21882 28376
rect 22094 28364 22100 28376
rect 22152 28364 22158 28416
rect 27065 28407 27123 28413
rect 27065 28373 27077 28407
rect 27111 28404 27123 28407
rect 27522 28404 27528 28416
rect 27111 28376 27528 28404
rect 27111 28373 27123 28376
rect 27065 28367 27123 28373
rect 27522 28364 27528 28376
rect 27580 28364 27586 28416
rect 27982 28404 27988 28416
rect 27943 28376 27988 28404
rect 27982 28364 27988 28376
rect 28040 28364 28046 28416
rect 30009 28407 30067 28413
rect 30009 28373 30021 28407
rect 30055 28404 30067 28407
rect 30374 28404 30380 28416
rect 30055 28376 30380 28404
rect 30055 28373 30067 28376
rect 30009 28367 30067 28373
rect 30374 28364 30380 28376
rect 30432 28364 30438 28416
rect 30650 28364 30656 28416
rect 30708 28404 30714 28416
rect 30761 28407 30819 28413
rect 30761 28404 30773 28407
rect 30708 28376 30773 28404
rect 30708 28364 30714 28376
rect 30761 28373 30773 28376
rect 30807 28373 30819 28407
rect 33226 28404 33232 28416
rect 33187 28376 33232 28404
rect 30761 28367 30819 28373
rect 33226 28364 33232 28376
rect 33284 28364 33290 28416
rect 34241 28407 34299 28413
rect 34241 28373 34253 28407
rect 34287 28404 34299 28407
rect 34974 28404 34980 28416
rect 34287 28376 34980 28404
rect 34287 28373 34299 28376
rect 34241 28367 34299 28373
rect 34974 28364 34980 28376
rect 35032 28364 35038 28416
rect 35342 28364 35348 28416
rect 35400 28404 35406 28416
rect 36265 28407 36323 28413
rect 36265 28404 36277 28407
rect 35400 28376 36277 28404
rect 35400 28364 35406 28376
rect 36265 28373 36277 28376
rect 36311 28373 36323 28407
rect 36265 28367 36323 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 10594 28160 10600 28212
rect 10652 28200 10658 28212
rect 23569 28203 23627 28209
rect 10652 28172 23520 28200
rect 10652 28160 10658 28172
rect 20162 28132 20168 28144
rect 17144 28104 19932 28132
rect 20123 28104 20168 28132
rect 17144 28076 17172 28104
rect 17126 28064 17132 28076
rect 17087 28036 17132 28064
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 17678 28064 17684 28076
rect 17512 28036 17684 28064
rect 17221 27999 17279 28005
rect 17221 27965 17233 27999
rect 17267 27965 17279 27999
rect 17221 27959 17279 27965
rect 16574 27820 16580 27872
rect 16632 27860 16638 27872
rect 17236 27860 17264 27959
rect 17512 27937 17540 28036
rect 17678 28024 17684 28036
rect 17736 28064 17742 28076
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 17736 28036 18521 28064
rect 17736 28024 17742 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 19705 28067 19763 28073
rect 19705 28033 19717 28067
rect 19751 28033 19763 28067
rect 19705 28027 19763 28033
rect 19797 28067 19855 28073
rect 19797 28033 19809 28067
rect 19843 28033 19855 28067
rect 19904 28064 19932 28104
rect 20162 28092 20168 28104
rect 20220 28092 20226 28144
rect 20548 28104 20852 28132
rect 20548 28064 20576 28104
rect 19904 28036 20576 28064
rect 19797 28027 19855 28033
rect 18414 27996 18420 28008
rect 18375 27968 18420 27996
rect 18414 27956 18420 27968
rect 18472 27956 18478 28008
rect 17497 27931 17555 27937
rect 17497 27897 17509 27931
rect 17543 27897 17555 27931
rect 17497 27891 17555 27897
rect 18877 27931 18935 27937
rect 18877 27897 18889 27931
rect 18923 27928 18935 27931
rect 19720 27928 19748 28027
rect 18923 27900 19748 27928
rect 18923 27897 18935 27900
rect 18877 27891 18935 27897
rect 17586 27860 17592 27872
rect 16632 27832 17592 27860
rect 16632 27820 16638 27832
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 19334 27820 19340 27872
rect 19392 27860 19398 27872
rect 19812 27860 19840 28027
rect 20622 28024 20628 28076
rect 20680 28064 20686 28076
rect 20824 28073 20852 28104
rect 23106 28092 23112 28144
rect 23164 28132 23170 28144
rect 23492 28132 23520 28172
rect 23569 28169 23581 28203
rect 23615 28200 23627 28203
rect 23658 28200 23664 28212
rect 23615 28172 23664 28200
rect 23615 28169 23627 28172
rect 23569 28163 23627 28169
rect 23658 28160 23664 28172
rect 23716 28160 23722 28212
rect 25774 28200 25780 28212
rect 25735 28172 25780 28200
rect 25774 28160 25780 28172
rect 25832 28160 25838 28212
rect 26145 28203 26203 28209
rect 26145 28169 26157 28203
rect 26191 28200 26203 28203
rect 26418 28200 26424 28212
rect 26191 28172 26424 28200
rect 26191 28169 26203 28172
rect 26145 28163 26203 28169
rect 26418 28160 26424 28172
rect 26476 28160 26482 28212
rect 27062 28160 27068 28212
rect 27120 28200 27126 28212
rect 27249 28203 27307 28209
rect 27249 28200 27261 28203
rect 27120 28172 27261 28200
rect 27120 28160 27126 28172
rect 27249 28169 27261 28172
rect 27295 28169 27307 28203
rect 27249 28163 27307 28169
rect 25038 28132 25044 28144
rect 23164 28104 23428 28132
rect 23492 28104 25044 28132
rect 23164 28092 23170 28104
rect 20809 28067 20867 28073
rect 20680 28036 20725 28064
rect 20680 28024 20686 28036
rect 20809 28033 20821 28067
rect 20855 28064 20867 28067
rect 21174 28064 21180 28076
rect 20855 28036 21180 28064
rect 20855 28033 20867 28036
rect 20809 28027 20867 28033
rect 21174 28024 21180 28036
rect 21232 28064 21238 28076
rect 23400 28073 23428 28104
rect 25038 28092 25044 28104
rect 25096 28132 25102 28144
rect 25096 28104 26004 28132
rect 25096 28092 25102 28104
rect 25976 28076 26004 28104
rect 21269 28067 21327 28073
rect 21269 28064 21281 28067
rect 21232 28036 21281 28064
rect 21232 28024 21238 28036
rect 21269 28033 21281 28036
rect 21315 28033 21327 28067
rect 21269 28027 21327 28033
rect 22465 28067 22523 28073
rect 22465 28033 22477 28067
rect 22511 28064 22523 28067
rect 23385 28067 23443 28073
rect 22511 28036 23336 28064
rect 22511 28033 22523 28036
rect 22465 28027 22523 28033
rect 20073 27999 20131 28005
rect 20073 27965 20085 27999
rect 20119 27996 20131 27999
rect 21450 27996 21456 28008
rect 20119 27968 21456 27996
rect 20119 27965 20131 27968
rect 20073 27959 20131 27965
rect 21450 27956 21456 27968
rect 21508 27956 21514 28008
rect 22646 27956 22652 28008
rect 22704 27996 22710 28008
rect 22741 27999 22799 28005
rect 22741 27996 22753 27999
rect 22704 27968 22753 27996
rect 22704 27956 22710 27968
rect 22741 27965 22753 27968
rect 22787 27996 22799 27999
rect 23201 27999 23259 28005
rect 23201 27996 23213 27999
rect 22787 27968 23213 27996
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 23201 27965 23213 27968
rect 23247 27965 23259 27999
rect 23308 27996 23336 28036
rect 23385 28033 23397 28067
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 24486 28024 24492 28076
rect 24544 28064 24550 28076
rect 24581 28067 24639 28073
rect 24581 28064 24593 28067
rect 24544 28036 24593 28064
rect 24544 28024 24550 28036
rect 24581 28033 24593 28036
rect 24627 28033 24639 28067
rect 25958 28064 25964 28076
rect 25871 28036 25964 28064
rect 24581 28027 24639 28033
rect 25958 28024 25964 28036
rect 26016 28024 26022 28076
rect 26237 28067 26295 28073
rect 26237 28033 26249 28067
rect 26283 28064 26295 28067
rect 26326 28064 26332 28076
rect 26283 28036 26332 28064
rect 26283 28033 26295 28036
rect 26237 28027 26295 28033
rect 26326 28024 26332 28036
rect 26384 28064 26390 28076
rect 27157 28067 27215 28073
rect 27157 28064 27169 28067
rect 26384 28036 27169 28064
rect 26384 28024 26390 28036
rect 27157 28033 27169 28036
rect 27203 28033 27215 28067
rect 27157 28027 27215 28033
rect 23566 27996 23572 28008
rect 23308 27968 23572 27996
rect 23201 27959 23259 27965
rect 23566 27956 23572 27968
rect 23624 27956 23630 28008
rect 24118 27956 24124 28008
rect 24176 27996 24182 28008
rect 24394 27996 24400 28008
rect 24176 27968 24400 27996
rect 24176 27956 24182 27968
rect 24394 27956 24400 27968
rect 24452 27956 24458 28008
rect 27264 27996 27292 28163
rect 28074 28160 28080 28212
rect 28132 28200 28138 28212
rect 28629 28203 28687 28209
rect 28629 28200 28641 28203
rect 28132 28172 28641 28200
rect 28132 28160 28138 28172
rect 28629 28169 28641 28172
rect 28675 28169 28687 28203
rect 28629 28163 28687 28169
rect 30561 28203 30619 28209
rect 30561 28169 30573 28203
rect 30607 28200 30619 28203
rect 30650 28200 30656 28212
rect 30607 28172 30656 28200
rect 30607 28169 30619 28172
rect 30561 28163 30619 28169
rect 30650 28160 30656 28172
rect 30708 28160 30714 28212
rect 30742 28160 30748 28212
rect 30800 28200 30806 28212
rect 31481 28203 31539 28209
rect 31481 28200 31493 28203
rect 30800 28172 31493 28200
rect 30800 28160 30806 28172
rect 31481 28169 31493 28172
rect 31527 28169 31539 28203
rect 31481 28163 31539 28169
rect 33689 28203 33747 28209
rect 33689 28169 33701 28203
rect 33735 28200 33747 28203
rect 34146 28200 34152 28212
rect 33735 28172 34152 28200
rect 33735 28169 33747 28172
rect 33689 28163 33747 28169
rect 34146 28160 34152 28172
rect 34204 28160 34210 28212
rect 34790 28200 34796 28212
rect 34751 28172 34796 28200
rect 34790 28160 34796 28172
rect 34848 28160 34854 28212
rect 35986 28200 35992 28212
rect 35947 28172 35992 28200
rect 35986 28160 35992 28172
rect 36044 28160 36050 28212
rect 27890 28092 27896 28144
rect 27948 28132 27954 28144
rect 28350 28132 28356 28144
rect 27948 28104 28120 28132
rect 28311 28104 28356 28132
rect 27948 28092 27954 28104
rect 27982 28064 27988 28076
rect 27943 28036 27988 28064
rect 27982 28024 27988 28036
rect 28040 28024 28046 28076
rect 28092 28073 28120 28104
rect 28350 28092 28356 28104
rect 28408 28092 28414 28144
rect 30285 28135 30343 28141
rect 30285 28101 30297 28135
rect 30331 28132 30343 28135
rect 30926 28132 30932 28144
rect 30331 28104 30932 28132
rect 30331 28101 30343 28104
rect 30285 28095 30343 28101
rect 30926 28092 30932 28104
rect 30984 28092 30990 28144
rect 32576 28135 32634 28141
rect 32576 28101 32588 28135
rect 32622 28132 32634 28135
rect 33226 28132 33232 28144
rect 32622 28104 33232 28132
rect 32622 28101 32634 28104
rect 32576 28095 32634 28101
rect 33226 28092 33232 28104
rect 33284 28092 33290 28144
rect 28078 28067 28136 28073
rect 28078 28033 28090 28067
rect 28124 28033 28136 28067
rect 28078 28027 28136 28033
rect 28258 28024 28264 28076
rect 28316 28064 28322 28076
rect 28316 28036 28409 28064
rect 28316 28024 28322 28036
rect 28442 28024 28448 28076
rect 28500 28073 28506 28076
rect 28500 28064 28508 28073
rect 29917 28067 29975 28073
rect 28500 28036 28545 28064
rect 28500 28027 28508 28036
rect 29917 28033 29929 28067
rect 29963 28033 29975 28067
rect 29917 28027 29975 28033
rect 28500 28024 28506 28027
rect 28276 27996 28304 28024
rect 27264 27968 28304 27996
rect 29932 27996 29960 28027
rect 30006 28024 30012 28076
rect 30064 28064 30070 28076
rect 30064 28036 30109 28064
rect 30064 28024 30070 28036
rect 30190 28024 30196 28076
rect 30248 28064 30254 28076
rect 30248 28036 30293 28064
rect 30248 28024 30254 28036
rect 30374 28024 30380 28076
rect 30432 28073 30438 28076
rect 30432 28064 30440 28073
rect 31018 28064 31024 28076
rect 30432 28036 30477 28064
rect 30979 28036 31024 28064
rect 30432 28027 30440 28036
rect 30432 28024 30438 28027
rect 31018 28024 31024 28036
rect 31076 28024 31082 28076
rect 34330 28064 34336 28076
rect 34291 28036 34336 28064
rect 34330 28024 34336 28036
rect 34388 28024 34394 28076
rect 34974 28064 34980 28076
rect 34935 28036 34980 28064
rect 34974 28024 34980 28036
rect 35032 28024 35038 28076
rect 36170 28064 36176 28076
rect 36131 28036 36176 28064
rect 36170 28024 36176 28036
rect 36228 28024 36234 28076
rect 36817 28067 36875 28073
rect 36817 28033 36829 28067
rect 36863 28064 36875 28067
rect 37550 28064 37556 28076
rect 36863 28036 37556 28064
rect 36863 28033 36875 28036
rect 36817 28027 36875 28033
rect 37550 28024 37556 28036
rect 37608 28024 37614 28076
rect 37642 28024 37648 28076
rect 37700 28064 37706 28076
rect 37700 28036 37745 28064
rect 37700 28024 37706 28036
rect 30466 27996 30472 28008
rect 29932 27968 30472 27996
rect 30466 27956 30472 27968
rect 30524 27956 30530 28008
rect 32030 27956 32036 28008
rect 32088 27996 32094 28008
rect 32309 27999 32367 28005
rect 32309 27996 32321 27999
rect 32088 27968 32321 27996
rect 32088 27956 32094 27968
rect 32309 27965 32321 27968
rect 32355 27965 32367 27999
rect 32309 27959 32367 27965
rect 37461 27999 37519 28005
rect 37461 27965 37473 27999
rect 37507 27996 37519 27999
rect 38010 27996 38016 28008
rect 37507 27968 38016 27996
rect 37507 27965 37519 27968
rect 37461 27959 37519 27965
rect 38010 27956 38016 27968
rect 38068 27956 38074 28008
rect 19981 27931 20039 27937
rect 19981 27897 19993 27931
rect 20027 27928 20039 27931
rect 20625 27931 20683 27937
rect 20625 27928 20637 27931
rect 20027 27900 20637 27928
rect 20027 27897 20039 27900
rect 19981 27891 20039 27897
rect 20625 27897 20637 27900
rect 20671 27897 20683 27931
rect 20625 27891 20683 27897
rect 21361 27931 21419 27937
rect 21361 27897 21373 27931
rect 21407 27928 21419 27931
rect 22094 27928 22100 27940
rect 21407 27900 22100 27928
rect 21407 27897 21419 27900
rect 21361 27891 21419 27897
rect 22094 27888 22100 27900
rect 22152 27928 22158 27940
rect 22554 27928 22560 27940
rect 22152 27900 22560 27928
rect 22152 27888 22158 27900
rect 22554 27888 22560 27900
rect 22612 27888 22618 27940
rect 24765 27931 24823 27937
rect 24765 27897 24777 27931
rect 24811 27928 24823 27931
rect 29178 27928 29184 27940
rect 24811 27900 29184 27928
rect 24811 27897 24823 27900
rect 24765 27891 24823 27897
rect 29178 27888 29184 27900
rect 29236 27888 29242 27940
rect 29270 27888 29276 27940
rect 29328 27928 29334 27940
rect 32214 27928 32220 27940
rect 29328 27900 32220 27928
rect 29328 27888 29334 27900
rect 32214 27888 32220 27900
rect 32272 27888 32278 27940
rect 34149 27931 34207 27937
rect 34149 27897 34161 27931
rect 34195 27928 34207 27931
rect 34606 27928 34612 27940
rect 34195 27900 34612 27928
rect 34195 27897 34207 27900
rect 34149 27891 34207 27897
rect 34606 27888 34612 27900
rect 34664 27888 34670 27940
rect 22278 27860 22284 27872
rect 19392 27832 19840 27860
rect 22239 27832 22284 27860
rect 19392 27820 19398 27832
rect 22278 27820 22284 27832
rect 22336 27820 22342 27872
rect 22649 27863 22707 27869
rect 22649 27829 22661 27863
rect 22695 27860 22707 27863
rect 23106 27860 23112 27872
rect 22695 27832 23112 27860
rect 22695 27829 22707 27832
rect 22649 27823 22707 27829
rect 23106 27820 23112 27832
rect 23164 27820 23170 27872
rect 25958 27820 25964 27872
rect 26016 27860 26022 27872
rect 29546 27860 29552 27872
rect 26016 27832 29552 27860
rect 26016 27820 26022 27832
rect 29546 27820 29552 27832
rect 29604 27820 29610 27872
rect 30926 27820 30932 27872
rect 30984 27860 30990 27872
rect 31113 27863 31171 27869
rect 31113 27860 31125 27863
rect 30984 27832 31125 27860
rect 30984 27820 30990 27832
rect 31113 27829 31125 27832
rect 31159 27829 31171 27863
rect 31113 27823 31171 27829
rect 36633 27863 36691 27869
rect 36633 27829 36645 27863
rect 36679 27860 36691 27863
rect 36722 27860 36728 27872
rect 36679 27832 36728 27860
rect 36679 27829 36691 27832
rect 36633 27823 36691 27829
rect 36722 27820 36728 27832
rect 36780 27820 36786 27872
rect 37458 27820 37464 27872
rect 37516 27860 37522 27872
rect 37829 27863 37887 27869
rect 37829 27860 37841 27863
rect 37516 27832 37841 27860
rect 37516 27820 37522 27832
rect 37829 27829 37841 27832
rect 37875 27829 37887 27863
rect 37829 27823 37887 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 18325 27659 18383 27665
rect 18325 27625 18337 27659
rect 18371 27656 18383 27659
rect 18414 27656 18420 27668
rect 18371 27628 18420 27656
rect 18371 27625 18383 27628
rect 18325 27619 18383 27625
rect 18414 27616 18420 27628
rect 18472 27616 18478 27668
rect 22646 27616 22652 27668
rect 22704 27656 22710 27668
rect 23109 27659 23167 27665
rect 23109 27656 23121 27659
rect 22704 27628 23121 27656
rect 22704 27616 22710 27628
rect 23109 27625 23121 27628
rect 23155 27625 23167 27659
rect 23109 27619 23167 27625
rect 27065 27659 27123 27665
rect 27065 27625 27077 27659
rect 27111 27656 27123 27659
rect 27246 27656 27252 27668
rect 27111 27628 27252 27656
rect 27111 27625 27123 27628
rect 27065 27619 27123 27625
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 34330 27656 34336 27668
rect 34291 27628 34336 27656
rect 34330 27616 34336 27628
rect 34388 27616 34394 27668
rect 35526 27616 35532 27668
rect 35584 27656 35590 27668
rect 35621 27659 35679 27665
rect 35621 27656 35633 27659
rect 35584 27628 35633 27656
rect 35584 27616 35590 27628
rect 35621 27625 35633 27628
rect 35667 27625 35679 27659
rect 36814 27656 36820 27668
rect 35621 27619 35679 27625
rect 36648 27628 36820 27656
rect 16853 27591 16911 27597
rect 16853 27557 16865 27591
rect 16899 27557 16911 27591
rect 17310 27588 17316 27600
rect 17271 27560 17316 27588
rect 16853 27551 16911 27557
rect 16574 27520 16580 27532
rect 16535 27492 16580 27520
rect 16574 27480 16580 27492
rect 16632 27480 16638 27532
rect 16868 27520 16896 27551
rect 17310 27548 17316 27560
rect 17368 27548 17374 27600
rect 17678 27588 17684 27600
rect 17639 27560 17684 27588
rect 17678 27548 17684 27560
rect 17736 27548 17742 27600
rect 18782 27548 18788 27600
rect 18840 27588 18846 27600
rect 20622 27588 20628 27600
rect 18840 27560 20628 27588
rect 18840 27548 18846 27560
rect 20622 27548 20628 27560
rect 20680 27548 20686 27600
rect 23566 27588 23572 27600
rect 23527 27560 23572 27588
rect 23566 27548 23572 27560
rect 23624 27548 23630 27600
rect 25682 27588 25688 27600
rect 25643 27560 25688 27588
rect 25682 27548 25688 27560
rect 25740 27548 25746 27600
rect 28534 27588 28540 27600
rect 26528 27560 28540 27588
rect 17589 27523 17647 27529
rect 17589 27520 17601 27523
rect 16868 27492 17601 27520
rect 17589 27489 17601 27492
rect 17635 27520 17647 27523
rect 17954 27520 17960 27532
rect 17635 27492 17960 27520
rect 17635 27489 17647 27492
rect 17589 27483 17647 27489
rect 17954 27480 17960 27492
rect 18012 27480 18018 27532
rect 23474 27480 23480 27532
rect 23532 27520 23538 27532
rect 23532 27492 23796 27520
rect 23532 27480 23538 27492
rect 16485 27455 16543 27461
rect 16485 27421 16497 27455
rect 16531 27421 16543 27455
rect 16485 27415 16543 27421
rect 17497 27455 17555 27461
rect 17497 27421 17509 27455
rect 17543 27452 17555 27455
rect 17678 27452 17684 27464
rect 17543 27424 17684 27452
rect 17543 27421 17555 27424
rect 17497 27415 17555 27421
rect 16500 27316 16528 27415
rect 17678 27412 17684 27424
rect 17736 27412 17742 27464
rect 17770 27412 17776 27464
rect 17828 27452 17834 27464
rect 18601 27455 18659 27461
rect 18601 27452 18613 27455
rect 17828 27424 17873 27452
rect 17972 27424 18613 27452
rect 17828 27412 17834 27424
rect 17586 27344 17592 27396
rect 17644 27384 17650 27396
rect 17972 27384 18000 27424
rect 18601 27421 18613 27424
rect 18647 27421 18659 27455
rect 18601 27415 18659 27421
rect 19978 27412 19984 27464
rect 20036 27452 20042 27464
rect 21729 27455 21787 27461
rect 21729 27452 21741 27455
rect 20036 27424 21741 27452
rect 20036 27412 20042 27424
rect 21729 27421 21741 27424
rect 21775 27421 21787 27455
rect 21729 27415 21787 27421
rect 21996 27455 22054 27461
rect 21996 27421 22008 27455
rect 22042 27452 22054 27455
rect 22278 27452 22284 27464
rect 22042 27424 22284 27452
rect 22042 27421 22054 27424
rect 21996 27415 22054 27421
rect 22278 27412 22284 27424
rect 22336 27412 22342 27464
rect 23569 27455 23627 27461
rect 23569 27421 23581 27455
rect 23615 27452 23627 27455
rect 23658 27452 23664 27464
rect 23615 27424 23664 27452
rect 23615 27421 23627 27424
rect 23569 27415 23627 27421
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 23768 27461 23796 27492
rect 24596 27492 26004 27520
rect 24596 27461 24624 27492
rect 23753 27455 23811 27461
rect 23753 27421 23765 27455
rect 23799 27421 23811 27455
rect 23753 27415 23811 27421
rect 24581 27455 24639 27461
rect 24581 27421 24593 27455
rect 24627 27421 24639 27455
rect 24581 27415 24639 27421
rect 24765 27455 24823 27461
rect 24765 27421 24777 27455
rect 24811 27452 24823 27455
rect 24946 27452 24952 27464
rect 24811 27424 24952 27452
rect 24811 27421 24823 27424
rect 24765 27415 24823 27421
rect 18322 27384 18328 27396
rect 17644 27356 18000 27384
rect 18283 27356 18328 27384
rect 17644 27344 17650 27356
rect 18322 27344 18328 27356
rect 18380 27344 18386 27396
rect 23768 27384 23796 27415
rect 24946 27412 24952 27424
rect 25004 27412 25010 27464
rect 25976 27461 26004 27492
rect 25961 27455 26019 27461
rect 25961 27421 25973 27455
rect 26007 27452 26019 27455
rect 26326 27452 26332 27464
rect 26007 27424 26332 27452
rect 26007 27421 26019 27424
rect 25961 27415 26019 27421
rect 26326 27412 26332 27424
rect 26384 27412 26390 27464
rect 26528 27461 26556 27560
rect 28534 27548 28540 27560
rect 28592 27548 28598 27600
rect 30006 27548 30012 27600
rect 30064 27588 30070 27600
rect 30466 27588 30472 27600
rect 30064 27560 30328 27588
rect 30427 27560 30472 27588
rect 30064 27548 30070 27560
rect 27338 27520 27344 27532
rect 26804 27492 27344 27520
rect 26804 27461 26832 27492
rect 27338 27480 27344 27492
rect 27396 27520 27402 27532
rect 27801 27523 27859 27529
rect 27801 27520 27813 27523
rect 27396 27492 27813 27520
rect 27396 27480 27402 27492
rect 27801 27489 27813 27492
rect 27847 27489 27859 27523
rect 27801 27483 27859 27489
rect 29638 27480 29644 27532
rect 29696 27520 29702 27532
rect 30101 27523 30159 27529
rect 30101 27520 30113 27523
rect 29696 27492 30113 27520
rect 29696 27480 29702 27492
rect 30101 27489 30113 27492
rect 30147 27520 30159 27523
rect 30190 27520 30196 27532
rect 30147 27492 30196 27520
rect 30147 27489 30159 27492
rect 30101 27483 30159 27489
rect 30190 27480 30196 27492
rect 30248 27480 30254 27532
rect 26513 27455 26571 27461
rect 26513 27421 26525 27455
rect 26559 27421 26571 27455
rect 26513 27415 26571 27421
rect 26789 27455 26847 27461
rect 26789 27421 26801 27455
rect 26835 27421 26847 27455
rect 26789 27415 26847 27421
rect 26881 27455 26939 27461
rect 26881 27421 26893 27455
rect 26927 27421 26939 27455
rect 27522 27452 27528 27464
rect 27483 27424 27528 27452
rect 26881 27415 26939 27421
rect 25222 27384 25228 27396
rect 23768 27356 25228 27384
rect 25222 27344 25228 27356
rect 25280 27344 25286 27396
rect 25685 27387 25743 27393
rect 25685 27353 25697 27387
rect 25731 27384 25743 27387
rect 26142 27384 26148 27396
rect 25731 27356 26148 27384
rect 25731 27353 25743 27356
rect 25685 27347 25743 27353
rect 26142 27344 26148 27356
rect 26200 27344 26206 27396
rect 26697 27387 26755 27393
rect 26697 27353 26709 27387
rect 26743 27353 26755 27387
rect 26896 27384 26924 27415
rect 27522 27412 27528 27424
rect 27580 27412 27586 27464
rect 27706 27452 27712 27464
rect 27667 27424 27712 27452
rect 27706 27412 27712 27424
rect 27764 27412 27770 27464
rect 27890 27412 27896 27464
rect 27948 27452 27954 27464
rect 28077 27455 28135 27461
rect 27948 27424 27993 27452
rect 27948 27412 27954 27424
rect 28077 27421 28089 27455
rect 28123 27452 28135 27455
rect 28166 27452 28172 27464
rect 28123 27424 28172 27452
rect 28123 27421 28135 27424
rect 28077 27415 28135 27421
rect 28166 27412 28172 27424
rect 28224 27412 28230 27464
rect 29178 27452 29184 27464
rect 29139 27424 29184 27452
rect 29178 27412 29184 27424
rect 29236 27412 29242 27464
rect 29730 27452 29736 27464
rect 29691 27424 29736 27452
rect 29730 27412 29736 27424
rect 29788 27412 29794 27464
rect 29914 27452 29920 27464
rect 29875 27424 29920 27452
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 30006 27412 30012 27464
rect 30064 27452 30070 27464
rect 30300 27461 30328 27560
rect 30466 27548 30472 27560
rect 30524 27548 30530 27600
rect 33318 27548 33324 27600
rect 33376 27588 33382 27600
rect 33413 27591 33471 27597
rect 33413 27588 33425 27591
rect 33376 27560 33425 27588
rect 33376 27548 33382 27560
rect 33413 27557 33425 27560
rect 33459 27588 33471 27591
rect 33686 27588 33692 27600
rect 33459 27560 33692 27588
rect 33459 27557 33471 27560
rect 33413 27551 33471 27557
rect 33686 27548 33692 27560
rect 33744 27548 33750 27600
rect 33594 27480 33600 27532
rect 33652 27520 33658 27532
rect 36648 27529 36676 27628
rect 36814 27616 36820 27628
rect 36872 27616 36878 27668
rect 36633 27523 36691 27529
rect 33652 27492 34192 27520
rect 33652 27480 33658 27492
rect 30285 27455 30343 27461
rect 30064 27424 30109 27452
rect 30064 27412 30070 27424
rect 30285 27421 30297 27455
rect 30331 27421 30343 27455
rect 30285 27415 30343 27421
rect 31205 27455 31263 27461
rect 31205 27421 31217 27455
rect 31251 27452 31263 27455
rect 32030 27452 32036 27464
rect 31251 27424 32036 27452
rect 31251 27421 31263 27424
rect 31205 27415 31263 27421
rect 32030 27412 32036 27424
rect 32088 27412 32094 27464
rect 34054 27452 34060 27464
rect 34015 27424 34060 27452
rect 34054 27412 34060 27424
rect 34112 27412 34118 27464
rect 34164 27461 34192 27492
rect 36633 27489 36645 27523
rect 36679 27489 36691 27523
rect 36633 27483 36691 27489
rect 34149 27455 34207 27461
rect 34149 27421 34161 27455
rect 34195 27421 34207 27455
rect 35066 27452 35072 27464
rect 35027 27424 35072 27452
rect 34149 27415 34207 27421
rect 35066 27412 35072 27424
rect 35124 27412 35130 27464
rect 35618 27452 35624 27464
rect 35579 27424 35624 27452
rect 35618 27412 35624 27424
rect 35676 27412 35682 27464
rect 35802 27452 35808 27464
rect 35763 27424 35808 27452
rect 35802 27412 35808 27424
rect 35860 27412 35866 27464
rect 36722 27412 36728 27464
rect 36780 27452 36786 27464
rect 36889 27455 36947 27461
rect 36889 27452 36901 27455
rect 36780 27424 36901 27452
rect 36780 27412 36786 27424
rect 36889 27421 36901 27424
rect 36935 27421 36947 27455
rect 36889 27415 36947 27421
rect 27724 27384 27752 27412
rect 31450 27387 31508 27393
rect 31450 27384 31462 27387
rect 26896 27356 27752 27384
rect 29012 27356 31462 27384
rect 26697 27347 26755 27353
rect 18506 27316 18512 27328
rect 16500 27288 18512 27316
rect 18506 27276 18512 27288
rect 18564 27276 18570 27328
rect 24670 27316 24676 27328
rect 24631 27288 24676 27316
rect 24670 27276 24676 27288
rect 24728 27276 24734 27328
rect 25869 27319 25927 27325
rect 25869 27285 25881 27319
rect 25915 27316 25927 27319
rect 26418 27316 26424 27328
rect 25915 27288 26424 27316
rect 25915 27285 25927 27288
rect 25869 27279 25927 27285
rect 26418 27276 26424 27288
rect 26476 27276 26482 27328
rect 26712 27316 26740 27347
rect 27430 27316 27436 27328
rect 26712 27288 27436 27316
rect 27430 27276 27436 27288
rect 27488 27276 27494 27328
rect 28166 27276 28172 27328
rect 28224 27316 28230 27328
rect 29012 27325 29040 27356
rect 31450 27353 31462 27356
rect 31496 27353 31508 27387
rect 33137 27387 33195 27393
rect 33137 27384 33149 27387
rect 31450 27347 31508 27353
rect 31726 27356 33149 27384
rect 28261 27319 28319 27325
rect 28261 27316 28273 27319
rect 28224 27288 28273 27316
rect 28224 27276 28230 27288
rect 28261 27285 28273 27288
rect 28307 27285 28319 27319
rect 28261 27279 28319 27285
rect 28997 27319 29055 27325
rect 28997 27285 29009 27319
rect 29043 27285 29055 27319
rect 28997 27279 29055 27285
rect 29086 27276 29092 27328
rect 29144 27316 29150 27328
rect 29454 27316 29460 27328
rect 29144 27288 29460 27316
rect 29144 27276 29150 27288
rect 29454 27276 29460 27288
rect 29512 27316 29518 27328
rect 30190 27316 30196 27328
rect 29512 27288 30196 27316
rect 29512 27276 29518 27288
rect 30190 27276 30196 27288
rect 30248 27276 30254 27328
rect 31294 27276 31300 27328
rect 31352 27316 31358 27328
rect 31726 27316 31754 27356
rect 33137 27353 33149 27356
rect 33183 27353 33195 27387
rect 33137 27347 33195 27353
rect 32582 27316 32588 27328
rect 31352 27288 31754 27316
rect 32543 27288 32588 27316
rect 31352 27276 31358 27288
rect 32582 27276 32588 27288
rect 32640 27276 32646 27328
rect 33152 27316 33180 27347
rect 34054 27316 34060 27328
rect 33152 27288 34060 27316
rect 34054 27276 34060 27288
rect 34112 27276 34118 27328
rect 34885 27319 34943 27325
rect 34885 27285 34897 27319
rect 34931 27316 34943 27319
rect 35342 27316 35348 27328
rect 34931 27288 35348 27316
rect 34931 27285 34943 27288
rect 34885 27279 34943 27285
rect 35342 27276 35348 27288
rect 35400 27276 35406 27328
rect 35989 27319 36047 27325
rect 35989 27285 36001 27319
rect 36035 27316 36047 27319
rect 36446 27316 36452 27328
rect 36035 27288 36452 27316
rect 36035 27285 36047 27288
rect 35989 27279 36047 27285
rect 36446 27276 36452 27288
rect 36504 27276 36510 27328
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 17313 27115 17371 27121
rect 17313 27081 17325 27115
rect 17359 27112 17371 27115
rect 17770 27112 17776 27124
rect 17359 27084 17776 27112
rect 17359 27081 17371 27084
rect 17313 27075 17371 27081
rect 17770 27072 17776 27084
rect 17828 27072 17834 27124
rect 22738 27112 22744 27124
rect 22699 27084 22744 27112
rect 22738 27072 22744 27084
rect 22796 27072 22802 27124
rect 25317 27115 25375 27121
rect 25317 27081 25329 27115
rect 25363 27112 25375 27115
rect 26326 27112 26332 27124
rect 26384 27121 26390 27124
rect 26384 27115 26403 27121
rect 25363 27084 26332 27112
rect 25363 27081 25375 27084
rect 25317 27075 25375 27081
rect 26326 27072 26332 27084
rect 26391 27081 26403 27115
rect 26384 27075 26403 27081
rect 27249 27115 27307 27121
rect 27249 27081 27261 27115
rect 27295 27112 27307 27115
rect 27430 27112 27436 27124
rect 27295 27084 27436 27112
rect 27295 27081 27307 27084
rect 27249 27075 27307 27081
rect 26384 27072 26390 27075
rect 27430 27072 27436 27084
rect 27488 27072 27494 27124
rect 28813 27115 28871 27121
rect 28813 27081 28825 27115
rect 28859 27112 28871 27115
rect 29730 27112 29736 27124
rect 28859 27084 29736 27112
rect 28859 27081 28871 27084
rect 28813 27075 28871 27081
rect 29730 27072 29736 27084
rect 29788 27072 29794 27124
rect 30282 27072 30288 27124
rect 30340 27072 30346 27124
rect 30374 27072 30380 27124
rect 30432 27112 30438 27124
rect 30469 27115 30527 27121
rect 30469 27112 30481 27115
rect 30432 27084 30481 27112
rect 30432 27072 30438 27084
rect 30469 27081 30481 27084
rect 30515 27112 30527 27115
rect 31018 27112 31024 27124
rect 30515 27084 31024 27112
rect 30515 27081 30527 27084
rect 30469 27075 30527 27081
rect 31018 27072 31024 27084
rect 31076 27072 31082 27124
rect 32214 27072 32220 27124
rect 32272 27112 32278 27124
rect 32585 27115 32643 27121
rect 32585 27112 32597 27115
rect 32272 27084 32597 27112
rect 32272 27072 32278 27084
rect 32585 27081 32597 27084
rect 32631 27112 32643 27115
rect 32766 27112 32772 27124
rect 32631 27084 32772 27112
rect 32631 27081 32643 27084
rect 32585 27075 32643 27081
rect 32766 27072 32772 27084
rect 32824 27072 32830 27124
rect 33873 27115 33931 27121
rect 33873 27081 33885 27115
rect 33919 27112 33931 27115
rect 35066 27112 35072 27124
rect 33919 27084 35072 27112
rect 33919 27081 33931 27084
rect 33873 27075 33931 27081
rect 35066 27072 35072 27084
rect 35124 27072 35130 27124
rect 35713 27115 35771 27121
rect 35713 27081 35725 27115
rect 35759 27112 35771 27115
rect 35802 27112 35808 27124
rect 35759 27084 35808 27112
rect 35759 27081 35771 27084
rect 35713 27075 35771 27081
rect 35802 27072 35808 27084
rect 35860 27112 35866 27124
rect 35860 27084 37504 27112
rect 35860 27072 35866 27084
rect 18601 27047 18659 27053
rect 18601 27013 18613 27047
rect 18647 27044 18659 27047
rect 19950 27047 20008 27053
rect 19950 27044 19962 27047
rect 18647 27016 19962 27044
rect 18647 27013 18659 27016
rect 18601 27007 18659 27013
rect 19950 27013 19962 27016
rect 19996 27013 20008 27047
rect 19950 27007 20008 27013
rect 24204 27047 24262 27053
rect 24204 27013 24216 27047
rect 24250 27044 24262 27047
rect 24670 27044 24676 27056
rect 24250 27016 24676 27044
rect 24250 27013 24262 27016
rect 24204 27007 24262 27013
rect 24670 27004 24676 27016
rect 24728 27004 24734 27056
rect 26142 27044 26148 27056
rect 26103 27016 26148 27044
rect 26142 27004 26148 27016
rect 26200 27004 26206 27056
rect 27890 27004 27896 27056
rect 27948 27044 27954 27056
rect 28445 27047 28503 27053
rect 28445 27044 28457 27047
rect 27948 27016 28457 27044
rect 27948 27004 27954 27016
rect 28445 27013 28457 27016
rect 28491 27013 28503 27047
rect 29914 27044 29920 27056
rect 28445 27007 28503 27013
rect 29196 27016 29920 27044
rect 17037 26979 17095 26985
rect 17037 26945 17049 26979
rect 17083 26976 17095 26979
rect 17126 26976 17132 26988
rect 17083 26948 17132 26976
rect 17083 26945 17095 26948
rect 17037 26939 17095 26945
rect 17126 26936 17132 26948
rect 17184 26936 17190 26988
rect 17954 26976 17960 26988
rect 17915 26948 17960 26976
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18506 26936 18512 26988
rect 18564 26976 18570 26988
rect 18877 26979 18935 26985
rect 18877 26976 18889 26979
rect 18564 26948 18889 26976
rect 18564 26936 18570 26948
rect 18877 26945 18889 26948
rect 18923 26945 18935 26979
rect 18877 26939 18935 26945
rect 18969 26979 19027 26985
rect 18969 26945 18981 26979
rect 19015 26945 19027 26979
rect 18969 26939 19027 26945
rect 17313 26911 17371 26917
rect 17313 26877 17325 26911
rect 17359 26908 17371 26911
rect 17494 26908 17500 26920
rect 17359 26880 17500 26908
rect 17359 26877 17371 26880
rect 17313 26871 17371 26877
rect 17494 26868 17500 26880
rect 17552 26868 17558 26920
rect 17770 26908 17776 26920
rect 17731 26880 17776 26908
rect 17770 26868 17776 26880
rect 17828 26868 17834 26920
rect 17129 26843 17187 26849
rect 17129 26809 17141 26843
rect 17175 26840 17187 26843
rect 18892 26840 18920 26939
rect 17175 26812 18920 26840
rect 18984 26840 19012 26939
rect 19058 26936 19064 26988
rect 19116 26976 19122 26988
rect 19116 26948 19161 26976
rect 19116 26936 19122 26948
rect 19242 26936 19248 26988
rect 19300 26976 19306 26988
rect 22005 26979 22063 26985
rect 19300 26948 19345 26976
rect 19444 26948 21128 26976
rect 19300 26936 19306 26948
rect 19334 26840 19340 26852
rect 18984 26812 19340 26840
rect 17175 26809 17187 26812
rect 17129 26803 17187 26809
rect 18141 26775 18199 26781
rect 18141 26741 18153 26775
rect 18187 26772 18199 26775
rect 18506 26772 18512 26784
rect 18187 26744 18512 26772
rect 18187 26741 18199 26744
rect 18141 26735 18199 26741
rect 18506 26732 18512 26744
rect 18564 26732 18570 26784
rect 18892 26772 18920 26812
rect 19334 26800 19340 26812
rect 19392 26800 19398 26852
rect 19444 26772 19472 26948
rect 19705 26911 19763 26917
rect 19705 26877 19717 26911
rect 19751 26877 19763 26911
rect 19705 26871 19763 26877
rect 18892 26744 19472 26772
rect 19720 26772 19748 26871
rect 21100 26784 21128 26948
rect 22005 26945 22017 26979
rect 22051 26945 22063 26979
rect 22186 26976 22192 26988
rect 22147 26948 22192 26976
rect 22005 26939 22063 26945
rect 22020 26908 22048 26939
rect 22186 26936 22192 26948
rect 22244 26936 22250 26988
rect 22554 26976 22560 26988
rect 22515 26948 22560 26976
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 26160 26976 26188 27004
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26160 26948 27169 26976
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 28166 26976 28172 26988
rect 28127 26948 28172 26976
rect 27157 26939 27215 26945
rect 28166 26936 28172 26948
rect 28224 26936 28230 26988
rect 28258 26936 28264 26988
rect 28316 26976 28322 26988
rect 28537 26979 28595 26985
rect 28316 26948 28361 26976
rect 28316 26936 28322 26948
rect 28537 26945 28549 26979
rect 28583 26945 28595 26979
rect 28537 26939 28595 26945
rect 28675 26979 28733 26985
rect 28675 26945 28687 26979
rect 28721 26976 28733 26979
rect 28994 26976 29000 26988
rect 28721 26948 29000 26976
rect 28721 26945 28733 26948
rect 28675 26939 28733 26945
rect 22094 26908 22100 26920
rect 22020 26880 22100 26908
rect 22094 26868 22100 26880
rect 22152 26868 22158 26920
rect 22281 26911 22339 26917
rect 22281 26877 22293 26911
rect 22327 26877 22339 26911
rect 22281 26871 22339 26877
rect 22373 26911 22431 26917
rect 22373 26877 22385 26911
rect 22419 26908 22431 26911
rect 22646 26908 22652 26920
rect 22419 26880 22652 26908
rect 22419 26877 22431 26880
rect 22373 26871 22431 26877
rect 21358 26800 21364 26852
rect 21416 26840 21422 26852
rect 22296 26840 22324 26871
rect 22646 26868 22652 26880
rect 22704 26868 22710 26920
rect 23937 26911 23995 26917
rect 23937 26877 23949 26911
rect 23983 26877 23995 26911
rect 23937 26871 23995 26877
rect 21416 26812 22324 26840
rect 21416 26800 21422 26812
rect 19978 26772 19984 26784
rect 19720 26744 19984 26772
rect 19978 26732 19984 26744
rect 20036 26732 20042 26784
rect 21082 26772 21088 26784
rect 21043 26744 21088 26772
rect 21082 26732 21088 26744
rect 21140 26732 21146 26784
rect 23952 26772 23980 26871
rect 27614 26868 27620 26920
rect 27672 26908 27678 26920
rect 28552 26908 28580 26939
rect 28994 26936 29000 26948
rect 29052 26976 29058 26988
rect 29196 26976 29224 27016
rect 29914 27004 29920 27016
rect 29972 27004 29978 27056
rect 30300 27044 30328 27072
rect 30300 27016 30604 27044
rect 29546 26976 29552 26988
rect 29052 26948 29224 26976
rect 29507 26948 29552 26976
rect 29052 26936 29058 26948
rect 29546 26936 29552 26948
rect 29604 26936 29610 26988
rect 30006 26976 30012 26988
rect 29656 26948 30012 26976
rect 29656 26908 29684 26948
rect 30006 26936 30012 26948
rect 30064 26936 30070 26988
rect 30190 26936 30196 26988
rect 30248 26976 30254 26988
rect 30576 26985 30604 27016
rect 31294 27004 31300 27056
rect 31352 27044 31358 27056
rect 31573 27047 31631 27053
rect 31573 27044 31585 27047
rect 31352 27016 31585 27044
rect 31352 27004 31358 27016
rect 31573 27013 31585 27016
rect 31619 27013 31631 27047
rect 31573 27007 31631 27013
rect 31757 27047 31815 27053
rect 31757 27013 31769 27047
rect 31803 27044 31815 27047
rect 32858 27044 32864 27056
rect 31803 27016 32864 27044
rect 31803 27013 31815 27016
rect 31757 27007 31815 27013
rect 32858 27004 32864 27016
rect 32916 27004 32922 27056
rect 36814 27044 36820 27056
rect 34348 27016 36820 27044
rect 30285 26979 30343 26985
rect 30285 26976 30297 26979
rect 30248 26948 30297 26976
rect 30248 26936 30254 26948
rect 30285 26945 30297 26948
rect 30331 26945 30343 26979
rect 30285 26939 30343 26945
rect 30561 26979 30619 26985
rect 30561 26945 30573 26979
rect 30607 26945 30619 26979
rect 32493 26979 32551 26985
rect 32493 26976 32505 26979
rect 30561 26939 30619 26945
rect 31726 26948 32505 26976
rect 27672 26880 29684 26908
rect 29825 26911 29883 26917
rect 27672 26868 27678 26880
rect 29825 26877 29837 26911
rect 29871 26908 29883 26911
rect 31726 26908 31754 26948
rect 32493 26945 32505 26948
rect 32539 26976 32551 26979
rect 33594 26976 33600 26988
rect 32539 26948 33600 26976
rect 32539 26945 32551 26948
rect 32493 26939 32551 26945
rect 33594 26936 33600 26948
rect 33652 26976 33658 26988
rect 34348 26985 34376 27016
rect 36814 27004 36820 27016
rect 36872 27004 36878 27056
rect 33689 26979 33747 26985
rect 33689 26976 33701 26979
rect 33652 26948 33701 26976
rect 33652 26936 33658 26948
rect 33689 26945 33701 26948
rect 33735 26945 33747 26979
rect 33689 26939 33747 26945
rect 34333 26979 34391 26985
rect 34333 26945 34345 26979
rect 34379 26945 34391 26979
rect 34333 26939 34391 26945
rect 34600 26979 34658 26985
rect 34600 26945 34612 26979
rect 34646 26976 34658 26979
rect 35342 26976 35348 26988
rect 34646 26948 35348 26976
rect 34646 26945 34658 26948
rect 34600 26939 34658 26945
rect 35342 26936 35348 26948
rect 35400 26936 35406 26988
rect 36354 26976 36360 26988
rect 36315 26948 36360 26976
rect 36354 26936 36360 26948
rect 36412 26936 36418 26988
rect 36446 26936 36452 26988
rect 36504 26976 36510 26988
rect 36630 26976 36636 26988
rect 36504 26948 36549 26976
rect 36591 26948 36636 26976
rect 36504 26936 36510 26948
rect 36630 26936 36636 26948
rect 36688 26936 36694 26988
rect 37476 26985 37504 27084
rect 37550 27072 37556 27124
rect 37608 27112 37614 27124
rect 37829 27115 37887 27121
rect 37829 27112 37841 27115
rect 37608 27084 37841 27112
rect 37608 27072 37614 27084
rect 37829 27081 37841 27084
rect 37875 27081 37887 27115
rect 37829 27075 37887 27081
rect 37461 26979 37519 26985
rect 37461 26945 37473 26979
rect 37507 26945 37519 26979
rect 37642 26976 37648 26988
rect 37603 26948 37648 26976
rect 37461 26939 37519 26945
rect 37642 26936 37648 26948
rect 37700 26936 37706 26988
rect 29871 26880 31754 26908
rect 33505 26911 33563 26917
rect 29871 26877 29883 26880
rect 29825 26871 29883 26877
rect 33505 26877 33517 26911
rect 33551 26877 33563 26911
rect 36372 26908 36400 26936
rect 38010 26908 38016 26920
rect 36372 26880 38016 26908
rect 33505 26871 33563 26877
rect 24670 26772 24676 26784
rect 23952 26744 24676 26772
rect 24670 26732 24676 26744
rect 24728 26732 24734 26784
rect 26329 26775 26387 26781
rect 26329 26741 26341 26775
rect 26375 26772 26387 26775
rect 26418 26772 26424 26784
rect 26375 26744 26424 26772
rect 26375 26741 26387 26744
rect 26329 26735 26387 26741
rect 26418 26732 26424 26744
rect 26476 26732 26482 26784
rect 26510 26732 26516 26784
rect 26568 26772 26574 26784
rect 26568 26744 26613 26772
rect 26568 26732 26574 26744
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 30285 26775 30343 26781
rect 30285 26772 30297 26775
rect 30156 26744 30297 26772
rect 30156 26732 30162 26744
rect 30285 26741 30297 26744
rect 30331 26741 30343 26775
rect 33520 26772 33548 26871
rect 38010 26868 38016 26880
rect 38068 26868 38074 26920
rect 36541 26843 36599 26849
rect 36541 26809 36553 26843
rect 36587 26840 36599 26843
rect 36906 26840 36912 26852
rect 36587 26812 36912 26840
rect 36587 26809 36599 26812
rect 36541 26803 36599 26809
rect 36906 26800 36912 26812
rect 36964 26800 36970 26852
rect 35526 26772 35532 26784
rect 33520 26744 35532 26772
rect 30285 26735 30343 26741
rect 35526 26732 35532 26744
rect 35584 26732 35590 26784
rect 36170 26772 36176 26784
rect 36131 26744 36176 26772
rect 36170 26732 36176 26744
rect 36228 26732 36234 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 17865 26571 17923 26577
rect 17865 26537 17877 26571
rect 17911 26568 17923 26571
rect 18322 26568 18328 26580
rect 17911 26540 18328 26568
rect 17911 26537 17923 26540
rect 17865 26531 17923 26537
rect 18322 26528 18328 26540
rect 18380 26568 18386 26580
rect 18601 26571 18659 26577
rect 18601 26568 18613 26571
rect 18380 26540 18613 26568
rect 18380 26528 18386 26540
rect 18601 26537 18613 26540
rect 18647 26537 18659 26571
rect 18601 26531 18659 26537
rect 18693 26571 18751 26577
rect 18693 26537 18705 26571
rect 18739 26568 18751 26571
rect 19058 26568 19064 26580
rect 18739 26540 19064 26568
rect 18739 26537 18751 26540
rect 18693 26531 18751 26537
rect 19058 26528 19064 26540
rect 19116 26528 19122 26580
rect 21358 26568 21364 26580
rect 21319 26540 21364 26568
rect 21358 26528 21364 26540
rect 21416 26528 21422 26580
rect 26142 26528 26148 26580
rect 26200 26568 26206 26580
rect 26513 26571 26571 26577
rect 26513 26568 26525 26571
rect 26200 26540 26525 26568
rect 26200 26528 26206 26540
rect 26513 26537 26525 26540
rect 26559 26537 26571 26571
rect 26513 26531 26571 26537
rect 27433 26571 27491 26577
rect 27433 26537 27445 26571
rect 27479 26568 27491 26571
rect 27706 26568 27712 26580
rect 27479 26540 27712 26568
rect 27479 26537 27491 26540
rect 27433 26531 27491 26537
rect 27706 26528 27712 26540
rect 27764 26528 27770 26580
rect 27890 26528 27896 26580
rect 27948 26568 27954 26580
rect 28077 26571 28135 26577
rect 28077 26568 28089 26571
rect 27948 26540 28089 26568
rect 27948 26528 27954 26540
rect 28077 26537 28089 26540
rect 28123 26537 28135 26571
rect 28994 26568 29000 26580
rect 28955 26540 29000 26568
rect 28077 26531 28135 26537
rect 28994 26528 29000 26540
rect 29052 26528 29058 26580
rect 36265 26571 36323 26577
rect 36265 26537 36277 26571
rect 36311 26568 36323 26571
rect 36354 26568 36360 26580
rect 36311 26540 36360 26568
rect 36311 26537 36323 26540
rect 36265 26531 36323 26537
rect 36354 26528 36360 26540
rect 36412 26528 36418 26580
rect 33318 26460 33324 26512
rect 33376 26500 33382 26512
rect 34606 26500 34612 26512
rect 33376 26472 34612 26500
rect 33376 26460 33382 26472
rect 34606 26460 34612 26472
rect 34664 26460 34670 26512
rect 36449 26503 36507 26509
rect 36449 26500 36461 26503
rect 35084 26472 36461 26500
rect 18230 26392 18236 26444
rect 18288 26432 18294 26444
rect 18782 26432 18788 26444
rect 18288 26404 18788 26432
rect 18288 26392 18294 26404
rect 18782 26392 18788 26404
rect 18840 26392 18846 26444
rect 30374 26432 30380 26444
rect 30335 26404 30380 26432
rect 30374 26392 30380 26404
rect 30432 26392 30438 26444
rect 32582 26392 32588 26444
rect 32640 26432 32646 26444
rect 33413 26435 33471 26441
rect 33413 26432 33425 26435
rect 32640 26404 33425 26432
rect 32640 26392 32646 26404
rect 33413 26401 33425 26404
rect 33459 26401 33471 26435
rect 33413 26395 33471 26401
rect 17865 26367 17923 26373
rect 17865 26333 17877 26367
rect 17911 26364 17923 26367
rect 17954 26364 17960 26376
rect 17911 26336 17960 26364
rect 17911 26333 17923 26336
rect 17865 26327 17923 26333
rect 17954 26324 17960 26336
rect 18012 26324 18018 26376
rect 18049 26367 18107 26373
rect 18049 26333 18061 26367
rect 18095 26333 18107 26367
rect 18506 26364 18512 26376
rect 18467 26336 18512 26364
rect 18049 26327 18107 26333
rect 17218 26256 17224 26308
rect 17276 26296 17282 26308
rect 17770 26296 17776 26308
rect 17276 26268 17776 26296
rect 17276 26256 17282 26268
rect 17770 26256 17776 26268
rect 17828 26296 17834 26308
rect 18064 26296 18092 26327
rect 18506 26324 18512 26336
rect 18564 26324 18570 26376
rect 21082 26324 21088 26376
rect 21140 26364 21146 26376
rect 21269 26367 21327 26373
rect 21269 26364 21281 26367
rect 21140 26336 21281 26364
rect 21140 26324 21146 26336
rect 21269 26333 21281 26336
rect 21315 26333 21327 26367
rect 21269 26327 21327 26333
rect 22925 26367 22983 26373
rect 22925 26333 22937 26367
rect 22971 26333 22983 26367
rect 23106 26364 23112 26376
rect 23067 26336 23112 26364
rect 22925 26327 22983 26333
rect 17828 26268 18092 26296
rect 17828 26256 17834 26268
rect 19242 26256 19248 26308
rect 19300 26296 19306 26308
rect 20070 26296 20076 26308
rect 19300 26268 20076 26296
rect 19300 26256 19306 26268
rect 20070 26256 20076 26268
rect 20128 26256 20134 26308
rect 22940 26296 22968 26327
rect 23106 26324 23112 26336
rect 23164 26324 23170 26376
rect 24670 26324 24676 26376
rect 24728 26364 24734 26376
rect 25133 26367 25191 26373
rect 25133 26364 25145 26367
rect 24728 26336 25145 26364
rect 24728 26324 24734 26336
rect 25133 26333 25145 26336
rect 25179 26364 25191 26367
rect 26234 26364 26240 26376
rect 25179 26336 26240 26364
rect 25179 26333 25191 26336
rect 25133 26327 25191 26333
rect 26234 26324 26240 26336
rect 26292 26324 26298 26376
rect 27154 26324 27160 26376
rect 27212 26364 27218 26376
rect 27341 26367 27399 26373
rect 27341 26364 27353 26367
rect 27212 26336 27353 26364
rect 27212 26324 27218 26336
rect 27341 26333 27353 26336
rect 27387 26333 27399 26367
rect 27341 26327 27399 26333
rect 27985 26367 28043 26373
rect 27985 26333 27997 26367
rect 28031 26364 28043 26367
rect 28534 26364 28540 26376
rect 28031 26336 28540 26364
rect 28031 26333 28043 26336
rect 27985 26327 28043 26333
rect 28534 26324 28540 26336
rect 28592 26324 28598 26376
rect 28905 26367 28963 26373
rect 28905 26333 28917 26367
rect 28951 26364 28963 26367
rect 28994 26364 29000 26376
rect 28951 26336 29000 26364
rect 28951 26333 28963 26336
rect 28905 26327 28963 26333
rect 28994 26324 29000 26336
rect 29052 26324 29058 26376
rect 30098 26364 30104 26376
rect 30059 26336 30104 26364
rect 30098 26324 30104 26336
rect 30156 26324 30162 26376
rect 30282 26364 30288 26376
rect 30243 26336 30288 26364
rect 30282 26324 30288 26336
rect 30340 26324 30346 26376
rect 33594 26364 33600 26376
rect 33555 26336 33600 26364
rect 33594 26324 33600 26336
rect 33652 26324 33658 26376
rect 35084 26373 35112 26472
rect 36449 26469 36461 26472
rect 36495 26469 36507 26503
rect 36449 26463 36507 26469
rect 38289 26503 38347 26509
rect 38289 26469 38301 26503
rect 38335 26469 38347 26503
rect 38289 26463 38347 26469
rect 35342 26432 35348 26444
rect 35176 26404 35348 26432
rect 35176 26373 35204 26404
rect 35342 26392 35348 26404
rect 35400 26392 35406 26444
rect 35529 26435 35587 26441
rect 35529 26401 35541 26435
rect 35575 26432 35587 26435
rect 36170 26432 36176 26444
rect 35575 26404 36176 26432
rect 35575 26401 35587 26404
rect 35529 26395 35587 26401
rect 36170 26392 36176 26404
rect 36228 26392 36234 26444
rect 36814 26392 36820 26444
rect 36872 26432 36878 26444
rect 36909 26435 36967 26441
rect 36909 26432 36921 26435
rect 36872 26404 36921 26432
rect 36872 26392 36878 26404
rect 36909 26401 36921 26404
rect 36955 26401 36967 26435
rect 36909 26395 36967 26401
rect 35069 26367 35127 26373
rect 35069 26333 35081 26367
rect 35115 26333 35127 26367
rect 35069 26327 35127 26333
rect 35161 26367 35219 26373
rect 35161 26333 35173 26367
rect 35207 26333 35219 26367
rect 35161 26327 35219 26333
rect 35250 26324 35256 26376
rect 35308 26364 35314 26376
rect 35618 26364 35624 26376
rect 35308 26336 35624 26364
rect 35308 26324 35314 26336
rect 35618 26324 35624 26336
rect 35676 26364 35682 26376
rect 38304 26364 38332 26463
rect 35676 26336 38332 26364
rect 35676 26324 35682 26336
rect 24486 26296 24492 26308
rect 22940 26268 24492 26296
rect 24486 26256 24492 26268
rect 24544 26256 24550 26308
rect 25400 26299 25458 26305
rect 25400 26265 25412 26299
rect 25446 26296 25458 26299
rect 25590 26296 25596 26308
rect 25446 26268 25596 26296
rect 25446 26265 25458 26268
rect 25400 26259 25458 26265
rect 25590 26256 25596 26268
rect 25648 26256 25654 26308
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26296 29975 26299
rect 30190 26296 30196 26308
rect 29963 26268 30196 26296
rect 29963 26265 29975 26268
rect 29917 26259 29975 26265
rect 30190 26256 30196 26268
rect 30248 26256 30254 26308
rect 31202 26296 31208 26308
rect 31163 26268 31208 26296
rect 31202 26256 31208 26268
rect 31260 26256 31266 26308
rect 33686 26256 33692 26308
rect 33744 26296 33750 26308
rect 33781 26299 33839 26305
rect 33781 26296 33793 26299
rect 33744 26268 33793 26296
rect 33744 26256 33750 26268
rect 33781 26265 33793 26268
rect 33827 26265 33839 26299
rect 33781 26259 33839 26265
rect 34606 26256 34612 26308
rect 34664 26296 34670 26308
rect 35371 26299 35429 26305
rect 35371 26296 35383 26299
rect 34664 26268 35383 26296
rect 34664 26256 34670 26268
rect 35371 26265 35383 26268
rect 35417 26265 35429 26299
rect 35371 26259 35429 26265
rect 35802 26256 35808 26308
rect 35860 26296 35866 26308
rect 36081 26299 36139 26305
rect 36081 26296 36093 26299
rect 35860 26268 36093 26296
rect 35860 26256 35866 26268
rect 36081 26265 36093 26268
rect 36127 26265 36139 26299
rect 36081 26259 36139 26265
rect 36170 26256 36176 26308
rect 36228 26296 36234 26308
rect 37154 26299 37212 26305
rect 37154 26296 37166 26299
rect 36228 26268 37166 26296
rect 36228 26256 36234 26268
rect 37154 26265 37166 26268
rect 37200 26265 37212 26299
rect 37154 26259 37212 26265
rect 22922 26188 22928 26240
rect 22980 26228 22986 26240
rect 23017 26231 23075 26237
rect 23017 26228 23029 26231
rect 22980 26200 23029 26228
rect 22980 26188 22986 26200
rect 23017 26197 23029 26200
rect 23063 26197 23075 26231
rect 23017 26191 23075 26197
rect 32030 26188 32036 26240
rect 32088 26228 32094 26240
rect 32493 26231 32551 26237
rect 32493 26228 32505 26231
rect 32088 26200 32505 26228
rect 32088 26188 32094 26200
rect 32493 26197 32505 26200
rect 32539 26197 32551 26231
rect 34882 26228 34888 26240
rect 34843 26200 34888 26228
rect 32493 26191 32551 26197
rect 34882 26188 34888 26200
rect 34940 26188 34946 26240
rect 36291 26231 36349 26237
rect 36291 26197 36303 26231
rect 36337 26228 36349 26231
rect 37274 26228 37280 26240
rect 36337 26200 37280 26228
rect 36337 26197 36349 26200
rect 36291 26191 36349 26197
rect 37274 26188 37280 26200
rect 37332 26188 37338 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 22925 26027 22983 26033
rect 22925 25993 22937 26027
rect 22971 26024 22983 26027
rect 23106 26024 23112 26036
rect 22971 25996 23112 26024
rect 22971 25993 22983 25996
rect 22925 25987 22983 25993
rect 23106 25984 23112 25996
rect 23164 25984 23170 26036
rect 24670 26024 24676 26036
rect 24631 25996 24676 26024
rect 24670 25984 24676 25996
rect 24728 25984 24734 26036
rect 25590 26024 25596 26036
rect 25551 25996 25596 26024
rect 25590 25984 25596 25996
rect 25648 25984 25654 26036
rect 29638 25984 29644 26036
rect 29696 26024 29702 26036
rect 34333 26027 34391 26033
rect 29696 25996 31754 26024
rect 29696 25984 29702 25996
rect 19334 25916 19340 25968
rect 19392 25956 19398 25968
rect 19392 25928 19840 25956
rect 19392 25916 19398 25928
rect 16942 25848 16948 25900
rect 17000 25888 17006 25900
rect 17589 25891 17647 25897
rect 17589 25888 17601 25891
rect 17000 25860 17601 25888
rect 17000 25848 17006 25860
rect 17589 25857 17601 25860
rect 17635 25888 17647 25891
rect 19702 25888 19708 25900
rect 17635 25860 19708 25888
rect 17635 25857 17647 25860
rect 17589 25851 17647 25857
rect 19702 25848 19708 25860
rect 19760 25848 19766 25900
rect 19812 25897 19840 25928
rect 22186 25916 22192 25968
rect 22244 25956 22250 25968
rect 22554 25956 22560 25968
rect 22244 25928 22560 25956
rect 22244 25916 22250 25928
rect 22554 25916 22560 25928
rect 22612 25916 22618 25968
rect 22773 25959 22831 25965
rect 22773 25925 22785 25959
rect 22819 25956 22831 25959
rect 26510 25956 26516 25968
rect 22819 25928 23152 25956
rect 22819 25925 22831 25928
rect 22773 25919 22831 25925
rect 23124 25900 23152 25928
rect 25608 25928 26516 25956
rect 19797 25891 19855 25897
rect 19797 25857 19809 25891
rect 19843 25857 19855 25891
rect 19797 25851 19855 25857
rect 19889 25891 19947 25897
rect 19889 25857 19901 25891
rect 19935 25857 19947 25891
rect 20070 25888 20076 25900
rect 20031 25860 20076 25888
rect 19889 25851 19947 25857
rect 17494 25820 17500 25832
rect 17455 25792 17500 25820
rect 17494 25780 17500 25792
rect 17552 25780 17558 25832
rect 19334 25780 19340 25832
rect 19392 25820 19398 25832
rect 19904 25820 19932 25851
rect 20070 25848 20076 25860
rect 20128 25848 20134 25900
rect 23106 25848 23112 25900
rect 23164 25848 23170 25900
rect 23382 25888 23388 25900
rect 23343 25860 23388 25888
rect 23382 25848 23388 25860
rect 23440 25848 23446 25900
rect 25608 25897 25636 25928
rect 26510 25916 26516 25928
rect 26568 25916 26574 25968
rect 30092 25959 30150 25965
rect 30092 25925 30104 25959
rect 30138 25956 30150 25959
rect 30190 25956 30196 25968
rect 30138 25928 30196 25956
rect 30138 25925 30150 25928
rect 30092 25919 30150 25925
rect 30190 25916 30196 25928
rect 30248 25916 30254 25968
rect 31726 25956 31754 25996
rect 34333 25993 34345 26027
rect 34379 26024 34391 26027
rect 34422 26024 34428 26036
rect 34379 25996 34428 26024
rect 34379 25993 34391 25996
rect 34333 25987 34391 25993
rect 34422 25984 34428 25996
rect 34480 26024 34486 26036
rect 36081 26027 36139 26033
rect 34480 25996 35894 26024
rect 34480 25984 34486 25996
rect 32401 25959 32459 25965
rect 32401 25956 32413 25959
rect 31726 25928 32413 25956
rect 32401 25925 32413 25928
rect 32447 25925 32459 25959
rect 34514 25956 34520 25968
rect 32401 25919 32459 25925
rect 32968 25928 34520 25956
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25682 25848 25688 25900
rect 25740 25888 25746 25900
rect 25740 25860 25785 25888
rect 25740 25848 25746 25860
rect 28810 25848 28816 25900
rect 28868 25888 28874 25900
rect 29089 25891 29147 25897
rect 29089 25888 29101 25891
rect 28868 25860 29101 25888
rect 28868 25848 28874 25860
rect 29089 25857 29101 25860
rect 29135 25888 29147 25891
rect 31386 25888 31392 25900
rect 29135 25860 31392 25888
rect 29135 25857 29147 25860
rect 29089 25851 29147 25857
rect 31386 25848 31392 25860
rect 31444 25888 31450 25900
rect 32968 25897 32996 25928
rect 34514 25916 34520 25928
rect 34572 25916 34578 25968
rect 34790 25916 34796 25968
rect 34848 25956 34854 25968
rect 35250 25956 35256 25968
rect 34848 25928 35256 25956
rect 34848 25916 34854 25928
rect 35250 25916 35256 25928
rect 35308 25916 35314 25968
rect 32309 25891 32367 25897
rect 32309 25888 32321 25891
rect 31444 25860 32321 25888
rect 31444 25848 31450 25860
rect 32309 25857 32321 25860
rect 32355 25857 32367 25891
rect 32309 25851 32367 25857
rect 32953 25891 33011 25897
rect 32953 25857 32965 25891
rect 32999 25857 33011 25891
rect 32953 25851 33011 25857
rect 33220 25891 33278 25897
rect 33220 25857 33232 25891
rect 33266 25888 33278 25891
rect 34882 25888 34888 25900
rect 33266 25860 34888 25888
rect 33266 25857 33278 25860
rect 33220 25851 33278 25857
rect 34882 25848 34888 25860
rect 34940 25848 34946 25900
rect 34977 25891 35035 25897
rect 34977 25857 34989 25891
rect 35023 25857 35035 25891
rect 34977 25851 35035 25857
rect 19392 25792 19932 25820
rect 19392 25780 19398 25792
rect 24394 25780 24400 25832
rect 24452 25820 24458 25832
rect 24946 25820 24952 25832
rect 24452 25792 24952 25820
rect 24452 25780 24458 25792
rect 24946 25780 24952 25792
rect 25004 25820 25010 25832
rect 25869 25823 25927 25829
rect 25869 25820 25881 25823
rect 25004 25792 25881 25820
rect 25004 25780 25010 25792
rect 25869 25789 25881 25792
rect 25915 25789 25927 25823
rect 25869 25783 25927 25789
rect 26326 25780 26332 25832
rect 26384 25820 26390 25832
rect 29362 25820 29368 25832
rect 26384 25792 29368 25820
rect 26384 25780 26390 25792
rect 29362 25780 29368 25792
rect 29420 25780 29426 25832
rect 29822 25820 29828 25832
rect 29783 25792 29828 25820
rect 29822 25780 29828 25792
rect 29880 25780 29886 25832
rect 34790 25820 34796 25832
rect 34751 25792 34796 25820
rect 34790 25780 34796 25792
rect 34848 25780 34854 25832
rect 17954 25752 17960 25764
rect 17915 25724 17960 25752
rect 17954 25712 17960 25724
rect 18012 25712 18018 25764
rect 31018 25712 31024 25764
rect 31076 25752 31082 25764
rect 31205 25755 31263 25761
rect 31205 25752 31217 25755
rect 31076 25724 31217 25752
rect 31076 25712 31082 25724
rect 31205 25721 31217 25724
rect 31251 25721 31263 25755
rect 34992 25752 35020 25851
rect 35866 25820 35894 25996
rect 36081 25993 36093 26027
rect 36127 26024 36139 26027
rect 36170 26024 36176 26036
rect 36127 25996 36176 26024
rect 36127 25993 36139 25996
rect 36081 25987 36139 25993
rect 36170 25984 36176 25996
rect 36228 25984 36234 26036
rect 37458 26024 37464 26036
rect 36280 25996 37464 26024
rect 36280 25897 36308 25996
rect 37458 25984 37464 25996
rect 37516 25984 37522 26036
rect 37829 25959 37887 25965
rect 37829 25956 37841 25959
rect 36924 25928 37841 25956
rect 36924 25897 36952 25928
rect 37829 25925 37841 25928
rect 37875 25925 37887 25959
rect 37829 25919 37887 25925
rect 36265 25891 36323 25897
rect 36265 25857 36277 25891
rect 36311 25857 36323 25891
rect 36265 25851 36323 25857
rect 36909 25891 36967 25897
rect 36909 25857 36921 25891
rect 36955 25857 36967 25891
rect 37642 25888 37648 25900
rect 37555 25860 37648 25888
rect 36909 25851 36967 25857
rect 37642 25848 37648 25860
rect 37700 25848 37706 25900
rect 36630 25820 36636 25832
rect 35866 25792 36636 25820
rect 36630 25780 36636 25792
rect 36688 25780 36694 25832
rect 37182 25780 37188 25832
rect 37240 25820 37246 25832
rect 37461 25823 37519 25829
rect 37461 25820 37473 25823
rect 37240 25792 37473 25820
rect 37240 25780 37246 25792
rect 37461 25789 37473 25792
rect 37507 25789 37519 25823
rect 37461 25783 37519 25789
rect 37660 25752 37688 25848
rect 34992 25724 37688 25752
rect 31205 25715 31263 25721
rect 19429 25687 19487 25693
rect 19429 25653 19441 25687
rect 19475 25684 19487 25687
rect 20070 25684 20076 25696
rect 19475 25656 20076 25684
rect 19475 25653 19487 25656
rect 19429 25647 19487 25653
rect 20070 25644 20076 25656
rect 20128 25644 20134 25696
rect 22741 25687 22799 25693
rect 22741 25653 22753 25687
rect 22787 25684 22799 25687
rect 23198 25684 23204 25696
rect 22787 25656 23204 25684
rect 22787 25653 22799 25656
rect 22741 25647 22799 25653
rect 23198 25644 23204 25656
rect 23256 25644 23262 25696
rect 29178 25684 29184 25696
rect 29139 25656 29184 25684
rect 29178 25644 29184 25656
rect 29236 25644 29242 25696
rect 29273 25687 29331 25693
rect 29273 25653 29285 25687
rect 29319 25684 29331 25687
rect 30742 25684 30748 25696
rect 29319 25656 30748 25684
rect 29319 25653 29331 25656
rect 29273 25647 29331 25653
rect 30742 25644 30748 25656
rect 30800 25644 30806 25696
rect 35161 25687 35219 25693
rect 35161 25653 35173 25687
rect 35207 25684 35219 25687
rect 35342 25684 35348 25696
rect 35207 25656 35348 25684
rect 35207 25653 35219 25656
rect 35161 25647 35219 25653
rect 35342 25644 35348 25656
rect 35400 25644 35406 25696
rect 36725 25687 36783 25693
rect 36725 25653 36737 25687
rect 36771 25684 36783 25687
rect 36998 25684 37004 25696
rect 36771 25656 37004 25684
rect 36771 25653 36783 25656
rect 36725 25647 36783 25653
rect 36998 25644 37004 25656
rect 37056 25644 37062 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 17218 25480 17224 25492
rect 17179 25452 17224 25480
rect 17218 25440 17224 25452
rect 17276 25440 17282 25492
rect 19702 25440 19708 25492
rect 19760 25480 19766 25492
rect 21177 25483 21235 25489
rect 21177 25480 21189 25483
rect 19760 25452 21189 25480
rect 19760 25440 19766 25452
rect 21177 25449 21189 25452
rect 21223 25449 21235 25483
rect 21177 25443 21235 25449
rect 21192 25412 21220 25443
rect 22094 25440 22100 25492
rect 22152 25480 22158 25492
rect 22189 25483 22247 25489
rect 22189 25480 22201 25483
rect 22152 25452 22201 25480
rect 22152 25440 22158 25452
rect 22189 25449 22201 25452
rect 22235 25449 22247 25483
rect 22189 25443 22247 25449
rect 22554 25440 22560 25492
rect 22612 25480 22618 25492
rect 22612 25452 24072 25480
rect 22612 25440 22618 25452
rect 22462 25412 22468 25424
rect 21192 25384 22468 25412
rect 22462 25372 22468 25384
rect 22520 25372 22526 25424
rect 17310 25304 17316 25356
rect 17368 25344 17374 25356
rect 17497 25347 17555 25353
rect 17497 25344 17509 25347
rect 17368 25316 17509 25344
rect 17368 25304 17374 25316
rect 17497 25313 17509 25316
rect 17543 25313 17555 25347
rect 17497 25307 17555 25313
rect 17589 25347 17647 25353
rect 17589 25313 17601 25347
rect 17635 25344 17647 25347
rect 17954 25344 17960 25356
rect 17635 25316 17960 25344
rect 17635 25313 17647 25316
rect 17589 25307 17647 25313
rect 17954 25304 17960 25316
rect 18012 25344 18018 25356
rect 18601 25347 18659 25353
rect 18601 25344 18613 25347
rect 18012 25316 18613 25344
rect 18012 25304 18018 25316
rect 18601 25313 18613 25316
rect 18647 25344 18659 25347
rect 19058 25344 19064 25356
rect 18647 25316 19064 25344
rect 18647 25313 18659 25316
rect 18601 25307 18659 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 21910 25344 21916 25356
rect 21652 25316 21916 25344
rect 17402 25276 17408 25288
rect 17363 25248 17408 25276
rect 17402 25236 17408 25248
rect 17460 25236 17466 25288
rect 17678 25236 17684 25288
rect 17736 25276 17742 25288
rect 18230 25276 18236 25288
rect 17736 25248 17781 25276
rect 18191 25248 18236 25276
rect 17736 25236 17742 25248
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 18693 25279 18751 25285
rect 18693 25245 18705 25279
rect 18739 25276 18751 25279
rect 18782 25276 18788 25288
rect 18739 25248 18788 25276
rect 18739 25245 18751 25248
rect 18693 25239 18751 25245
rect 18782 25236 18788 25248
rect 18840 25236 18846 25288
rect 19797 25279 19855 25285
rect 19797 25245 19809 25279
rect 19843 25276 19855 25279
rect 19886 25276 19892 25288
rect 19843 25248 19892 25276
rect 19843 25245 19855 25248
rect 19797 25239 19855 25245
rect 19886 25236 19892 25248
rect 19944 25236 19950 25288
rect 20070 25285 20076 25288
rect 20064 25276 20076 25285
rect 20031 25248 20076 25276
rect 20064 25239 20076 25248
rect 20070 25236 20076 25239
rect 20128 25236 20134 25288
rect 21652 25285 21680 25316
rect 21910 25304 21916 25316
rect 21968 25304 21974 25356
rect 22572 25344 22600 25440
rect 24044 25421 24072 25452
rect 24486 25440 24492 25492
rect 24544 25480 24550 25492
rect 25501 25483 25559 25489
rect 25501 25480 25513 25483
rect 24544 25452 25513 25480
rect 24544 25440 24550 25452
rect 25501 25449 25513 25452
rect 25547 25449 25559 25483
rect 27154 25480 27160 25492
rect 27115 25452 27160 25480
rect 25501 25443 25559 25449
rect 27154 25440 27160 25452
rect 27212 25440 27218 25492
rect 28994 25480 29000 25492
rect 28955 25452 29000 25480
rect 28994 25440 29000 25452
rect 29052 25480 29058 25492
rect 29270 25480 29276 25492
rect 29052 25452 29276 25480
rect 29052 25440 29058 25452
rect 29270 25440 29276 25452
rect 29328 25440 29334 25492
rect 29362 25440 29368 25492
rect 29420 25480 29426 25492
rect 31386 25480 31392 25492
rect 29420 25452 31248 25480
rect 31347 25452 31392 25480
rect 29420 25440 29426 25452
rect 24029 25415 24087 25421
rect 24029 25381 24041 25415
rect 24075 25381 24087 25415
rect 24029 25375 24087 25381
rect 22020 25316 22600 25344
rect 24044 25344 24072 25375
rect 24578 25372 24584 25424
rect 24636 25412 24642 25424
rect 24765 25415 24823 25421
rect 24765 25412 24777 25415
rect 24636 25384 24777 25412
rect 24636 25372 24642 25384
rect 24765 25381 24777 25384
rect 24811 25381 24823 25415
rect 26326 25412 26332 25424
rect 24765 25375 24823 25381
rect 25608 25384 26332 25412
rect 24044 25316 24808 25344
rect 21637 25279 21695 25285
rect 21637 25245 21649 25279
rect 21683 25245 21695 25279
rect 21818 25276 21824 25288
rect 21779 25248 21824 25276
rect 21637 25239 21695 25245
rect 21818 25236 21824 25248
rect 21876 25236 21882 25288
rect 22020 25285 22048 25316
rect 22005 25279 22063 25285
rect 22005 25245 22017 25279
rect 22051 25245 22063 25279
rect 22646 25276 22652 25288
rect 22607 25248 22652 25276
rect 22005 25239 22063 25245
rect 22646 25236 22652 25248
rect 22704 25236 22710 25288
rect 22922 25285 22928 25288
rect 22916 25276 22928 25285
rect 22883 25248 22928 25276
rect 22916 25239 22928 25248
rect 22922 25236 22928 25239
rect 22980 25236 22986 25288
rect 23198 25236 23204 25288
rect 23256 25276 23262 25288
rect 24486 25276 24492 25288
rect 23256 25248 24492 25276
rect 23256 25236 23262 25248
rect 24486 25236 24492 25248
rect 24544 25276 24550 25288
rect 24581 25279 24639 25285
rect 24581 25276 24593 25279
rect 24544 25248 24593 25276
rect 24544 25236 24550 25248
rect 24581 25245 24593 25248
rect 24627 25245 24639 25279
rect 24581 25239 24639 25245
rect 24673 25279 24731 25285
rect 24673 25245 24685 25279
rect 24719 25245 24731 25279
rect 24780 25276 24808 25316
rect 24854 25304 24860 25356
rect 24912 25344 24918 25356
rect 25608 25353 25636 25384
rect 26326 25372 26332 25384
rect 26384 25372 26390 25424
rect 25593 25347 25651 25353
rect 25593 25344 25605 25347
rect 24912 25316 25605 25344
rect 24912 25304 24918 25316
rect 25593 25313 25605 25316
rect 25639 25313 25651 25347
rect 25593 25307 25651 25313
rect 26145 25347 26203 25353
rect 26145 25313 26157 25347
rect 26191 25344 26203 25347
rect 26234 25344 26240 25356
rect 26191 25316 26240 25344
rect 26191 25313 26203 25316
rect 26145 25307 26203 25313
rect 26234 25304 26240 25316
rect 26292 25344 26298 25356
rect 27172 25344 27200 25440
rect 27341 25415 27399 25421
rect 27341 25381 27353 25415
rect 27387 25381 27399 25415
rect 31220 25412 31248 25452
rect 31386 25440 31392 25452
rect 31444 25440 31450 25492
rect 33318 25480 33324 25492
rect 31726 25452 33324 25480
rect 31726 25412 31754 25452
rect 33318 25440 33324 25452
rect 33376 25440 33382 25492
rect 33502 25440 33508 25492
rect 33560 25480 33566 25492
rect 34054 25480 34060 25492
rect 33560 25452 34060 25480
rect 33560 25440 33566 25452
rect 34054 25440 34060 25452
rect 34112 25440 34118 25492
rect 31220 25384 31754 25412
rect 27341 25375 27399 25381
rect 26292 25316 27200 25344
rect 27356 25344 27384 25375
rect 27356 25316 28028 25344
rect 26292 25304 26298 25316
rect 25317 25279 25375 25285
rect 25317 25276 25329 25279
rect 24780 25248 25329 25276
rect 24673 25239 24731 25245
rect 25317 25245 25329 25248
rect 25363 25245 25375 25279
rect 25317 25239 25375 25245
rect 25409 25279 25467 25285
rect 25409 25245 25421 25279
rect 25455 25245 25467 25279
rect 25409 25239 25467 25245
rect 18248 25208 18276 25236
rect 19242 25208 19248 25220
rect 18248 25180 19248 25208
rect 19242 25168 19248 25180
rect 19300 25168 19306 25220
rect 21358 25168 21364 25220
rect 21416 25208 21422 25220
rect 21913 25211 21971 25217
rect 21913 25208 21925 25211
rect 21416 25180 21925 25208
rect 21416 25168 21422 25180
rect 21913 25177 21925 25180
rect 21959 25177 21971 25211
rect 21913 25171 21971 25177
rect 23106 25168 23112 25220
rect 23164 25208 23170 25220
rect 24688 25208 24716 25239
rect 23164 25180 24716 25208
rect 23164 25168 23170 25180
rect 24762 25168 24768 25220
rect 24820 25208 24826 25220
rect 25424 25208 25452 25239
rect 25866 25236 25872 25288
rect 25924 25276 25930 25288
rect 26329 25279 26387 25285
rect 26329 25276 26341 25279
rect 25924 25248 26341 25276
rect 25924 25236 25930 25248
rect 26329 25245 26341 25248
rect 26375 25276 26387 25279
rect 26510 25276 26516 25288
rect 26375 25248 26516 25276
rect 26375 25245 26387 25248
rect 26329 25239 26387 25245
rect 26510 25236 26516 25248
rect 26568 25236 26574 25288
rect 27798 25276 27804 25288
rect 27759 25248 27804 25276
rect 27798 25236 27804 25248
rect 27856 25236 27862 25288
rect 28000 25285 28028 25316
rect 28994 25304 29000 25356
rect 29052 25344 29058 25356
rect 29822 25344 29828 25356
rect 29052 25316 29828 25344
rect 29052 25304 29058 25316
rect 29822 25304 29828 25316
rect 29880 25344 29886 25356
rect 30009 25347 30067 25353
rect 30009 25344 30021 25347
rect 29880 25316 30021 25344
rect 29880 25304 29886 25316
rect 30009 25313 30021 25316
rect 30055 25313 30067 25347
rect 30009 25307 30067 25313
rect 33796 25316 34560 25344
rect 27985 25279 28043 25285
rect 27985 25245 27997 25279
rect 28031 25245 28043 25279
rect 27985 25239 28043 25245
rect 32033 25279 32091 25285
rect 32033 25245 32045 25279
rect 32079 25276 32091 25279
rect 33796 25276 33824 25316
rect 34532 25288 34560 25316
rect 36722 25304 36728 25356
rect 36780 25344 36786 25356
rect 36909 25347 36967 25353
rect 36909 25344 36921 25347
rect 36780 25316 36921 25344
rect 36780 25304 36786 25316
rect 36909 25313 36921 25316
rect 36955 25313 36967 25347
rect 36909 25307 36967 25313
rect 32079 25248 33824 25276
rect 33873 25279 33931 25285
rect 32079 25245 32091 25248
rect 32033 25239 32091 25245
rect 33873 25245 33885 25279
rect 33919 25245 33931 25279
rect 33873 25239 33931 25245
rect 24820 25180 25452 25208
rect 26528 25208 26556 25236
rect 26973 25211 27031 25217
rect 26528 25180 26648 25208
rect 24820 25168 24826 25180
rect 18598 25100 18604 25152
rect 18656 25140 18662 25152
rect 18877 25143 18935 25149
rect 18877 25140 18889 25143
rect 18656 25112 18889 25140
rect 18656 25100 18662 25112
rect 18877 25109 18889 25112
rect 18923 25109 18935 25143
rect 18877 25103 18935 25109
rect 22002 25100 22008 25152
rect 22060 25140 22066 25152
rect 22278 25140 22284 25152
rect 22060 25112 22284 25140
rect 22060 25100 22066 25112
rect 22278 25100 22284 25112
rect 22336 25100 22342 25152
rect 26510 25140 26516 25152
rect 26471 25112 26516 25140
rect 26510 25100 26516 25112
rect 26568 25100 26574 25152
rect 26620 25140 26648 25180
rect 26973 25177 26985 25211
rect 27019 25208 27031 25211
rect 27614 25208 27620 25220
rect 27019 25180 27620 25208
rect 27019 25177 27031 25180
rect 26973 25171 27031 25177
rect 27614 25168 27620 25180
rect 27672 25168 27678 25220
rect 27173 25143 27231 25149
rect 27173 25140 27185 25143
rect 26620 25112 27185 25140
rect 27173 25109 27185 25112
rect 27219 25109 27231 25143
rect 27890 25140 27896 25152
rect 27851 25112 27896 25140
rect 27173 25103 27231 25109
rect 27890 25100 27896 25112
rect 27948 25100 27954 25152
rect 28000 25140 28028 25239
rect 28810 25208 28816 25220
rect 28771 25180 28816 25208
rect 28810 25168 28816 25180
rect 28868 25168 28874 25220
rect 29029 25211 29087 25217
rect 29029 25208 29041 25211
rect 29028 25177 29041 25208
rect 29075 25208 29087 25211
rect 29362 25208 29368 25220
rect 29075 25180 29368 25208
rect 29075 25177 29087 25180
rect 29028 25171 29087 25177
rect 29028 25140 29056 25171
rect 29362 25168 29368 25180
rect 29420 25168 29426 25220
rect 30276 25211 30334 25217
rect 30276 25177 30288 25211
rect 30322 25208 30334 25211
rect 30834 25208 30840 25220
rect 30322 25180 30840 25208
rect 30322 25177 30334 25180
rect 30276 25171 30334 25177
rect 30834 25168 30840 25180
rect 30892 25168 30898 25220
rect 32300 25211 32358 25217
rect 32300 25177 32312 25211
rect 32346 25208 32358 25211
rect 32950 25208 32956 25220
rect 32346 25180 32956 25208
rect 32346 25177 32358 25180
rect 32300 25171 32358 25177
rect 32950 25168 32956 25180
rect 33008 25168 33014 25220
rect 33318 25168 33324 25220
rect 33376 25208 33382 25220
rect 33888 25208 33916 25239
rect 34514 25236 34520 25288
rect 34572 25276 34578 25288
rect 34885 25279 34943 25285
rect 34885 25276 34897 25279
rect 34572 25248 34897 25276
rect 34572 25236 34578 25248
rect 34885 25245 34897 25248
rect 34931 25276 34943 25279
rect 36170 25276 36176 25288
rect 34931 25248 36176 25276
rect 34931 25245 34943 25248
rect 34885 25239 34943 25245
rect 36170 25236 36176 25248
rect 36228 25276 36234 25288
rect 36740 25276 36768 25304
rect 36228 25248 36768 25276
rect 36228 25236 36234 25248
rect 36998 25236 37004 25288
rect 37056 25276 37062 25288
rect 37165 25279 37223 25285
rect 37165 25276 37177 25279
rect 37056 25248 37177 25276
rect 37056 25236 37062 25248
rect 37165 25245 37177 25248
rect 37211 25245 37223 25279
rect 37165 25239 37223 25245
rect 33376 25180 33916 25208
rect 33376 25168 33382 25180
rect 34974 25168 34980 25220
rect 35032 25208 35038 25220
rect 35130 25211 35188 25217
rect 35130 25208 35142 25211
rect 35032 25180 35142 25208
rect 35032 25168 35038 25180
rect 35130 25177 35142 25180
rect 35176 25177 35188 25211
rect 35130 25171 35188 25177
rect 28000 25112 29056 25140
rect 29181 25143 29239 25149
rect 29181 25109 29193 25143
rect 29227 25140 29239 25143
rect 30006 25140 30012 25152
rect 29227 25112 30012 25140
rect 29227 25109 29239 25112
rect 29181 25103 29239 25109
rect 30006 25100 30012 25112
rect 30064 25100 30070 25152
rect 33413 25143 33471 25149
rect 33413 25109 33425 25143
rect 33459 25140 33471 25143
rect 33870 25140 33876 25152
rect 33459 25112 33876 25140
rect 33459 25109 33471 25112
rect 33413 25103 33471 25109
rect 33870 25100 33876 25112
rect 33928 25100 33934 25152
rect 36265 25143 36323 25149
rect 36265 25109 36277 25143
rect 36311 25140 36323 25143
rect 37182 25140 37188 25152
rect 36311 25112 37188 25140
rect 36311 25109 36323 25112
rect 36265 25103 36323 25109
rect 37182 25100 37188 25112
rect 37240 25100 37246 25152
rect 37642 25100 37648 25152
rect 37700 25140 37706 25152
rect 38289 25143 38347 25149
rect 38289 25140 38301 25143
rect 37700 25112 38301 25140
rect 37700 25100 37706 25112
rect 38289 25109 38301 25112
rect 38335 25109 38347 25143
rect 38289 25103 38347 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 16960 24908 18000 24936
rect 16117 24803 16175 24809
rect 16117 24769 16129 24803
rect 16163 24769 16175 24803
rect 16298 24800 16304 24812
rect 16259 24772 16304 24800
rect 16117 24763 16175 24769
rect 16132 24664 16160 24763
rect 16298 24760 16304 24772
rect 16356 24800 16362 24812
rect 16960 24800 16988 24908
rect 17402 24868 17408 24880
rect 17052 24840 17408 24868
rect 17052 24809 17080 24840
rect 17402 24828 17408 24840
rect 17460 24868 17466 24880
rect 17862 24868 17868 24880
rect 17460 24840 17868 24868
rect 17460 24828 17466 24840
rect 17862 24828 17868 24840
rect 17920 24828 17926 24880
rect 16356 24772 16988 24800
rect 17037 24803 17095 24809
rect 16356 24760 16362 24772
rect 17037 24769 17049 24803
rect 17083 24769 17095 24803
rect 17770 24800 17776 24812
rect 17731 24772 17776 24800
rect 17037 24763 17095 24769
rect 17770 24760 17776 24772
rect 17828 24760 17834 24812
rect 17972 24809 18000 24908
rect 22002 24896 22008 24948
rect 22060 24936 22066 24948
rect 22060 24908 22232 24936
rect 22060 24896 22066 24908
rect 22204 24877 22232 24908
rect 24486 24896 24492 24948
rect 24544 24936 24550 24948
rect 24857 24939 24915 24945
rect 24857 24936 24869 24939
rect 24544 24908 24869 24936
rect 24544 24896 24550 24908
rect 24857 24905 24869 24908
rect 24903 24905 24915 24939
rect 24857 24899 24915 24905
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 28534 24936 28540 24948
rect 27672 24908 28540 24936
rect 27672 24896 27678 24908
rect 28534 24896 28540 24908
rect 28592 24896 28598 24948
rect 34885 24939 34943 24945
rect 34885 24905 34897 24939
rect 34931 24936 34943 24939
rect 34974 24936 34980 24948
rect 34931 24908 34980 24936
rect 34931 24905 34943 24908
rect 34885 24899 34943 24905
rect 34974 24896 34980 24908
rect 35032 24896 35038 24948
rect 37182 24896 37188 24948
rect 37240 24936 37246 24948
rect 37645 24939 37703 24945
rect 37645 24936 37657 24939
rect 37240 24908 37657 24936
rect 37240 24896 37246 24908
rect 37645 24905 37657 24908
rect 37691 24905 37703 24939
rect 37645 24899 37703 24905
rect 22189 24871 22247 24877
rect 22189 24837 22201 24871
rect 22235 24868 22247 24871
rect 22925 24871 22983 24877
rect 22925 24868 22937 24871
rect 22235 24840 22937 24868
rect 22235 24837 22247 24840
rect 22189 24831 22247 24837
rect 22925 24837 22937 24840
rect 22971 24837 22983 24871
rect 24670 24868 24676 24880
rect 22925 24831 22983 24837
rect 23492 24840 24676 24868
rect 17957 24803 18015 24809
rect 17957 24769 17969 24803
rect 18003 24769 18015 24803
rect 18598 24800 18604 24812
rect 18559 24772 18604 24800
rect 17957 24763 18015 24769
rect 18598 24760 18604 24772
rect 18656 24760 18662 24812
rect 18782 24760 18788 24812
rect 18840 24800 18846 24812
rect 18877 24803 18935 24809
rect 18877 24800 18889 24803
rect 18840 24772 18889 24800
rect 18840 24760 18846 24772
rect 18877 24769 18889 24772
rect 18923 24769 18935 24803
rect 19058 24800 19064 24812
rect 19019 24772 19064 24800
rect 18877 24763 18935 24769
rect 19058 24760 19064 24772
rect 19116 24760 19122 24812
rect 19978 24800 19984 24812
rect 19904 24772 19984 24800
rect 16209 24735 16267 24741
rect 16209 24701 16221 24735
rect 16255 24732 16267 24735
rect 17313 24735 17371 24741
rect 17313 24732 17325 24735
rect 16255 24704 17325 24732
rect 16255 24701 16267 24704
rect 16209 24695 16267 24701
rect 17313 24701 17325 24704
rect 17359 24732 17371 24735
rect 18690 24732 18696 24744
rect 17359 24704 18696 24732
rect 17359 24701 17371 24704
rect 17313 24695 17371 24701
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 17034 24664 17040 24676
rect 16132 24636 17040 24664
rect 17034 24624 17040 24636
rect 17092 24624 17098 24676
rect 17221 24667 17279 24673
rect 17221 24633 17233 24667
rect 17267 24664 17279 24667
rect 18800 24664 18828 24760
rect 19904 24741 19932 24772
rect 19978 24760 19984 24772
rect 20036 24760 20042 24812
rect 20162 24809 20168 24812
rect 20156 24763 20168 24809
rect 20220 24800 20226 24812
rect 22005 24803 22063 24809
rect 20220 24772 20256 24800
rect 20162 24760 20168 24763
rect 20220 24760 20226 24772
rect 22005 24769 22017 24803
rect 22051 24800 22063 24803
rect 22094 24800 22100 24812
rect 22051 24772 22100 24800
rect 22051 24769 22063 24772
rect 22005 24763 22063 24769
rect 22094 24760 22100 24772
rect 22152 24760 22158 24812
rect 22462 24760 22468 24812
rect 22520 24800 22526 24812
rect 23492 24809 23520 24840
rect 24670 24828 24676 24840
rect 24728 24828 24734 24880
rect 26510 24868 26516 24880
rect 25884 24840 26516 24868
rect 22833 24803 22891 24809
rect 22833 24800 22845 24803
rect 22520 24772 22845 24800
rect 22520 24760 22526 24772
rect 22833 24769 22845 24772
rect 22879 24769 22891 24803
rect 22833 24763 22891 24769
rect 23477 24803 23535 24809
rect 23477 24769 23489 24803
rect 23523 24769 23535 24803
rect 23477 24763 23535 24769
rect 23744 24803 23802 24809
rect 23744 24769 23756 24803
rect 23790 24800 23802 24803
rect 24486 24800 24492 24812
rect 23790 24772 24492 24800
rect 23790 24769 23802 24772
rect 23744 24763 23802 24769
rect 24486 24760 24492 24772
rect 24544 24760 24550 24812
rect 25317 24803 25375 24809
rect 25317 24769 25329 24803
rect 25363 24769 25375 24803
rect 25317 24763 25375 24769
rect 25501 24803 25559 24809
rect 25501 24769 25513 24803
rect 25547 24800 25559 24803
rect 25884 24800 25912 24840
rect 26510 24828 26516 24840
rect 26568 24828 26574 24880
rect 33870 24868 33876 24880
rect 33152 24840 33876 24868
rect 25547 24772 25912 24800
rect 25547 24769 25559 24772
rect 25501 24763 25559 24769
rect 19889 24735 19947 24741
rect 19889 24701 19901 24735
rect 19935 24701 19947 24735
rect 19889 24695 19947 24701
rect 17267 24636 18828 24664
rect 18877 24667 18935 24673
rect 17267 24633 17279 24636
rect 17221 24627 17279 24633
rect 18877 24633 18889 24667
rect 18923 24664 18935 24667
rect 19334 24664 19340 24676
rect 18923 24636 19340 24664
rect 18923 24633 18935 24636
rect 18877 24627 18935 24633
rect 19334 24624 19340 24636
rect 19392 24624 19398 24676
rect 17129 24599 17187 24605
rect 17129 24565 17141 24599
rect 17175 24596 17187 24599
rect 17310 24596 17316 24608
rect 17175 24568 17316 24596
rect 17175 24565 17187 24568
rect 17129 24559 17187 24565
rect 17310 24556 17316 24568
rect 17368 24556 17374 24608
rect 18141 24599 18199 24605
rect 18141 24565 18153 24599
rect 18187 24596 18199 24599
rect 18782 24596 18788 24608
rect 18187 24568 18788 24596
rect 18187 24565 18199 24568
rect 18141 24559 18199 24565
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 19904 24596 19932 24695
rect 21818 24692 21824 24744
rect 21876 24732 21882 24744
rect 22373 24735 22431 24741
rect 22373 24732 22385 24735
rect 21876 24704 22385 24732
rect 21876 24692 21882 24704
rect 22373 24701 22385 24704
rect 22419 24701 22431 24735
rect 22373 24695 22431 24701
rect 22646 24664 22652 24676
rect 20824 24636 22652 24664
rect 20824 24596 20852 24636
rect 22646 24624 22652 24636
rect 22704 24624 22710 24676
rect 25332 24664 25360 24763
rect 25958 24760 25964 24812
rect 26016 24800 26022 24812
rect 26016 24772 26061 24800
rect 26016 24760 26022 24772
rect 26418 24760 26424 24812
rect 26476 24800 26482 24812
rect 27157 24803 27215 24809
rect 27157 24800 27169 24803
rect 26476 24772 27169 24800
rect 26476 24760 26482 24772
rect 27157 24769 27169 24772
rect 27203 24769 27215 24803
rect 27157 24763 27215 24769
rect 27424 24803 27482 24809
rect 27424 24769 27436 24803
rect 27470 24800 27482 24803
rect 27890 24800 27896 24812
rect 27470 24772 27896 24800
rect 27470 24769 27482 24772
rect 27424 24763 27482 24769
rect 27890 24760 27896 24772
rect 27948 24760 27954 24812
rect 28534 24760 28540 24812
rect 28592 24800 28598 24812
rect 29253 24803 29311 24809
rect 29253 24800 29265 24803
rect 28592 24772 29265 24800
rect 28592 24760 28598 24772
rect 29253 24769 29265 24772
rect 29299 24769 29311 24803
rect 29253 24763 29311 24769
rect 30742 24760 30748 24812
rect 30800 24800 30806 24812
rect 30837 24803 30895 24809
rect 30837 24800 30849 24803
rect 30800 24772 30849 24800
rect 30800 24760 30806 24772
rect 30837 24769 30849 24772
rect 30883 24769 30895 24803
rect 30837 24763 30895 24769
rect 31021 24803 31079 24809
rect 31021 24769 31033 24803
rect 31067 24769 31079 24803
rect 31021 24763 31079 24769
rect 31665 24803 31723 24809
rect 31665 24769 31677 24803
rect 31711 24800 31723 24803
rect 32306 24800 32312 24812
rect 31711 24772 32312 24800
rect 31711 24769 31723 24772
rect 31665 24763 31723 24769
rect 26237 24735 26295 24741
rect 26237 24701 26249 24735
rect 26283 24732 26295 24735
rect 26326 24732 26332 24744
rect 26283 24704 26332 24732
rect 26283 24701 26295 24704
rect 26237 24695 26295 24701
rect 26326 24692 26332 24704
rect 26384 24692 26390 24744
rect 28994 24692 29000 24744
rect 29052 24732 29058 24744
rect 29052 24704 29097 24732
rect 29052 24692 29058 24704
rect 30006 24692 30012 24744
rect 30064 24732 30070 24744
rect 30282 24732 30288 24744
rect 30064 24704 30288 24732
rect 30064 24692 30070 24704
rect 30282 24692 30288 24704
rect 30340 24732 30346 24744
rect 31036 24732 31064 24763
rect 32306 24760 32312 24772
rect 32364 24760 32370 24812
rect 32585 24803 32643 24809
rect 32585 24769 32597 24803
rect 32631 24769 32643 24803
rect 32585 24763 32643 24769
rect 32861 24803 32919 24809
rect 32861 24769 32873 24803
rect 32907 24800 32919 24803
rect 33152 24800 33180 24840
rect 33870 24828 33876 24840
rect 33928 24828 33934 24880
rect 37829 24871 37887 24877
rect 37829 24868 37841 24871
rect 36648 24840 37841 24868
rect 33686 24800 33692 24812
rect 32907 24772 33180 24800
rect 33647 24772 33692 24800
rect 32907 24769 32919 24772
rect 32861 24763 32919 24769
rect 30340 24704 31064 24732
rect 30340 24692 30346 24704
rect 31938 24692 31944 24744
rect 31996 24732 32002 24744
rect 32600 24732 32628 24763
rect 33686 24760 33692 24772
rect 33744 24760 33750 24812
rect 35069 24803 35127 24809
rect 35069 24769 35081 24803
rect 35115 24800 35127 24803
rect 35342 24800 35348 24812
rect 35115 24772 35348 24800
rect 35115 24769 35127 24772
rect 35069 24763 35127 24769
rect 35342 24760 35348 24772
rect 35400 24760 35406 24812
rect 36449 24803 36507 24809
rect 36449 24769 36461 24803
rect 36495 24800 36507 24803
rect 36648 24800 36676 24840
rect 37829 24837 37841 24840
rect 37875 24868 37887 24871
rect 38286 24868 38292 24880
rect 37875 24840 38292 24868
rect 37875 24837 37887 24840
rect 37829 24831 37887 24837
rect 38286 24828 38292 24840
rect 38344 24828 38350 24880
rect 36495 24772 36676 24800
rect 36725 24803 36783 24809
rect 36495 24769 36507 24772
rect 36449 24763 36507 24769
rect 36725 24769 36737 24803
rect 36771 24800 36783 24803
rect 37458 24800 37464 24812
rect 36771 24772 37464 24800
rect 36771 24769 36783 24772
rect 36725 24763 36783 24769
rect 37458 24760 37464 24772
rect 37516 24800 37522 24812
rect 37642 24800 37648 24812
rect 37516 24772 37648 24800
rect 37516 24760 37522 24772
rect 37642 24760 37648 24772
rect 37700 24760 37706 24812
rect 37737 24803 37795 24809
rect 37737 24769 37749 24803
rect 37783 24769 37795 24803
rect 37737 24763 37795 24769
rect 31996 24704 32628 24732
rect 32769 24735 32827 24741
rect 31996 24692 32002 24704
rect 32769 24701 32781 24735
rect 32815 24732 32827 24735
rect 33410 24732 33416 24744
rect 32815 24704 33416 24732
rect 32815 24701 32827 24704
rect 32769 24695 32827 24701
rect 33410 24692 33416 24704
rect 33468 24692 33474 24744
rect 36633 24735 36691 24741
rect 36633 24701 36645 24735
rect 36679 24732 36691 24735
rect 37550 24732 37556 24744
rect 36679 24704 37556 24732
rect 36679 24701 36691 24704
rect 36633 24695 36691 24701
rect 37550 24692 37556 24704
rect 37608 24732 37614 24744
rect 37752 24732 37780 24763
rect 37608 24704 37780 24732
rect 37608 24692 37614 24704
rect 26145 24667 26203 24673
rect 26145 24664 26157 24667
rect 25332 24636 26157 24664
rect 26145 24633 26157 24636
rect 26191 24633 26203 24667
rect 30834 24664 30840 24676
rect 30795 24636 30840 24664
rect 26145 24627 26203 24633
rect 30834 24624 30840 24636
rect 30892 24624 30898 24676
rect 32950 24624 32956 24676
rect 33008 24664 33014 24676
rect 33505 24667 33563 24673
rect 33505 24664 33517 24667
rect 33008 24636 33517 24664
rect 33008 24624 33014 24636
rect 33505 24633 33517 24636
rect 33551 24633 33563 24667
rect 36906 24664 36912 24676
rect 36867 24636 36912 24664
rect 33505 24627 33563 24633
rect 36906 24624 36912 24636
rect 36964 24624 36970 24676
rect 37274 24624 37280 24676
rect 37332 24664 37338 24676
rect 38013 24667 38071 24673
rect 38013 24664 38025 24667
rect 37332 24636 38025 24664
rect 37332 24624 37338 24636
rect 38013 24633 38025 24636
rect 38059 24633 38071 24667
rect 38013 24627 38071 24633
rect 21266 24596 21272 24608
rect 19904 24568 20852 24596
rect 21227 24568 21272 24596
rect 21266 24556 21272 24568
rect 21324 24556 21330 24608
rect 25317 24599 25375 24605
rect 25317 24565 25329 24599
rect 25363 24596 25375 24599
rect 25406 24596 25412 24608
rect 25363 24568 25412 24596
rect 25363 24565 25375 24568
rect 25317 24559 25375 24565
rect 25406 24556 25412 24568
rect 25464 24556 25470 24608
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 26053 24599 26111 24605
rect 26053 24596 26065 24599
rect 25924 24568 26065 24596
rect 25924 24556 25930 24568
rect 26053 24565 26065 24568
rect 26099 24565 26111 24599
rect 26053 24559 26111 24565
rect 29270 24556 29276 24608
rect 29328 24596 29334 24608
rect 30377 24599 30435 24605
rect 30377 24596 30389 24599
rect 29328 24568 30389 24596
rect 29328 24556 29334 24568
rect 30377 24565 30389 24568
rect 30423 24565 30435 24599
rect 30377 24559 30435 24565
rect 31481 24599 31539 24605
rect 31481 24565 31493 24599
rect 31527 24596 31539 24599
rect 32122 24596 32128 24608
rect 31527 24568 32128 24596
rect 31527 24565 31539 24568
rect 31481 24559 31539 24565
rect 32122 24556 32128 24568
rect 32180 24556 32186 24608
rect 32582 24596 32588 24608
rect 32543 24568 32588 24596
rect 32582 24556 32588 24568
rect 32640 24556 32646 24608
rect 33042 24596 33048 24608
rect 33003 24568 33048 24596
rect 33042 24556 33048 24568
rect 33100 24556 33106 24608
rect 36725 24599 36783 24605
rect 36725 24565 36737 24599
rect 36771 24596 36783 24599
rect 37182 24596 37188 24608
rect 36771 24568 37188 24596
rect 36771 24565 36783 24568
rect 36725 24559 36783 24565
rect 37182 24556 37188 24568
rect 37240 24556 37246 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 16298 24352 16304 24404
rect 16356 24392 16362 24404
rect 17037 24395 17095 24401
rect 17037 24392 17049 24395
rect 16356 24364 17049 24392
rect 16356 24352 16362 24364
rect 17037 24361 17049 24364
rect 17083 24361 17095 24395
rect 17037 24355 17095 24361
rect 17129 24395 17187 24401
rect 17129 24361 17141 24395
rect 17175 24392 17187 24395
rect 17678 24392 17684 24404
rect 17175 24364 17684 24392
rect 17175 24361 17187 24364
rect 17129 24355 17187 24361
rect 16942 24188 16948 24200
rect 16903 24160 16948 24188
rect 16942 24148 16948 24160
rect 17000 24148 17006 24200
rect 17052 24120 17080 24355
rect 17678 24352 17684 24364
rect 17736 24352 17742 24404
rect 19521 24395 19579 24401
rect 19521 24361 19533 24395
rect 19567 24392 19579 24395
rect 20162 24392 20168 24404
rect 19567 24364 20168 24392
rect 19567 24361 19579 24364
rect 19521 24355 19579 24361
rect 20162 24352 20168 24364
rect 20220 24352 20226 24404
rect 22278 24392 22284 24404
rect 22239 24364 22284 24392
rect 22278 24352 22284 24364
rect 22336 24352 22342 24404
rect 24486 24352 24492 24404
rect 24544 24392 24550 24404
rect 24581 24395 24639 24401
rect 24581 24392 24593 24395
rect 24544 24364 24593 24392
rect 24544 24352 24550 24364
rect 24581 24361 24593 24364
rect 24627 24361 24639 24395
rect 24581 24355 24639 24361
rect 26234 24352 26240 24404
rect 26292 24352 26298 24404
rect 26510 24352 26516 24404
rect 26568 24392 26574 24404
rect 27249 24395 27307 24401
rect 27249 24392 27261 24395
rect 26568 24364 27261 24392
rect 26568 24352 26574 24364
rect 27249 24361 27261 24364
rect 27295 24361 27307 24395
rect 27249 24355 27307 24361
rect 27341 24395 27399 24401
rect 27341 24361 27353 24395
rect 27387 24392 27399 24395
rect 27798 24392 27804 24404
rect 27387 24364 27804 24392
rect 27387 24361 27399 24364
rect 27341 24355 27399 24361
rect 27798 24352 27804 24364
rect 27856 24352 27862 24404
rect 28534 24392 28540 24404
rect 28495 24364 28540 24392
rect 28534 24352 28540 24364
rect 28592 24352 28598 24404
rect 28905 24395 28963 24401
rect 28905 24361 28917 24395
rect 28951 24392 28963 24395
rect 28951 24364 29132 24392
rect 28951 24361 28963 24364
rect 28905 24355 28963 24361
rect 17310 24284 17316 24336
rect 17368 24324 17374 24336
rect 18785 24327 18843 24333
rect 18785 24324 18797 24327
rect 17368 24296 18797 24324
rect 17368 24284 17374 24296
rect 17218 24256 17224 24268
rect 17179 24228 17224 24256
rect 17218 24216 17224 24228
rect 17276 24256 17282 24268
rect 17494 24256 17500 24268
rect 17276 24228 17500 24256
rect 17276 24216 17282 24228
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17972 24265 18000 24296
rect 18785 24293 18797 24296
rect 18831 24293 18843 24327
rect 23750 24324 23756 24336
rect 23711 24296 23756 24324
rect 18785 24287 18843 24293
rect 23750 24284 23756 24296
rect 23808 24284 23814 24336
rect 26252 24324 26280 24352
rect 26697 24327 26755 24333
rect 26697 24324 26709 24327
rect 26252 24296 26709 24324
rect 26697 24293 26709 24296
rect 26743 24293 26755 24327
rect 29104 24324 29132 24364
rect 29178 24352 29184 24404
rect 29236 24392 29242 24404
rect 30101 24395 30159 24401
rect 30101 24392 30113 24395
rect 29236 24364 30113 24392
rect 29236 24352 29242 24364
rect 30101 24361 30113 24364
rect 30147 24361 30159 24395
rect 33410 24392 33416 24404
rect 33371 24364 33416 24392
rect 30101 24355 30159 24361
rect 33410 24352 33416 24364
rect 33468 24352 33474 24404
rect 37550 24392 37556 24404
rect 37511 24364 37556 24392
rect 37550 24352 37556 24364
rect 37608 24352 37614 24404
rect 29362 24324 29368 24336
rect 29104 24296 29368 24324
rect 26697 24287 26755 24293
rect 29362 24284 29368 24296
rect 29420 24324 29426 24336
rect 29420 24296 29960 24324
rect 29420 24284 29426 24296
rect 17957 24259 18015 24265
rect 17957 24225 17969 24259
rect 18003 24225 18015 24259
rect 17957 24219 18015 24225
rect 19426 24216 19432 24268
rect 19484 24256 19490 24268
rect 21085 24259 21143 24265
rect 19484 24228 19932 24256
rect 19484 24216 19490 24228
rect 17862 24188 17868 24200
rect 17823 24160 17868 24188
rect 17862 24148 17868 24160
rect 17920 24148 17926 24200
rect 18690 24188 18696 24200
rect 18651 24160 18696 24188
rect 18690 24148 18696 24160
rect 18748 24148 18754 24200
rect 18782 24148 18788 24200
rect 18840 24188 18846 24200
rect 19904 24197 19932 24228
rect 21085 24225 21097 24259
rect 21131 24256 21143 24259
rect 22554 24256 22560 24268
rect 21131 24228 22560 24256
rect 21131 24225 21143 24228
rect 21085 24219 21143 24225
rect 18877 24191 18935 24197
rect 18877 24188 18889 24191
rect 18840 24160 18889 24188
rect 18840 24148 18846 24160
rect 18877 24157 18889 24160
rect 18923 24157 18935 24191
rect 18877 24151 18935 24157
rect 19797 24191 19855 24197
rect 19797 24157 19809 24191
rect 19843 24157 19855 24191
rect 19797 24151 19855 24157
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24157 19947 24191
rect 19889 24151 19947 24157
rect 19812 24120 19840 24151
rect 19978 24148 19984 24200
rect 20036 24188 20042 24200
rect 20165 24191 20223 24197
rect 20036 24160 20081 24188
rect 20036 24148 20042 24160
rect 20165 24157 20177 24191
rect 20211 24188 20223 24191
rect 20254 24188 20260 24200
rect 20211 24160 20260 24188
rect 20211 24157 20223 24160
rect 20165 24151 20223 24157
rect 20254 24148 20260 24160
rect 20312 24148 20318 24200
rect 20993 24191 21051 24197
rect 20993 24157 21005 24191
rect 21039 24188 21051 24191
rect 21266 24188 21272 24200
rect 21039 24160 21272 24188
rect 21039 24157 21051 24160
rect 20993 24151 21051 24157
rect 21008 24120 21036 24151
rect 21266 24148 21272 24160
rect 21324 24148 21330 24200
rect 21634 24188 21640 24200
rect 21595 24160 21640 24188
rect 21634 24148 21640 24160
rect 21692 24148 21698 24200
rect 21745 24197 21773 24228
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 22925 24259 22983 24265
rect 22925 24225 22937 24259
rect 22971 24256 22983 24259
rect 23198 24256 23204 24268
rect 22971 24228 23204 24256
rect 22971 24225 22983 24228
rect 22925 24219 22983 24225
rect 21730 24191 21788 24197
rect 21730 24157 21742 24191
rect 21776 24157 21788 24191
rect 22002 24188 22008 24200
rect 21963 24160 22008 24188
rect 21730 24151 21788 24157
rect 22002 24148 22008 24160
rect 22060 24148 22066 24200
rect 22094 24148 22100 24200
rect 22152 24197 22158 24200
rect 22152 24191 22201 24197
rect 22152 24157 22155 24191
rect 22189 24188 22201 24191
rect 22940 24188 22968 24219
rect 23198 24216 23204 24228
rect 23256 24216 23262 24268
rect 23566 24216 23572 24268
rect 23624 24256 23630 24268
rect 23624 24228 24072 24256
rect 23624 24216 23630 24228
rect 23106 24188 23112 24200
rect 22189 24160 22968 24188
rect 23067 24160 23112 24188
rect 22189 24157 22201 24160
rect 22152 24151 22201 24157
rect 22152 24148 22158 24151
rect 23106 24148 23112 24160
rect 23164 24148 23170 24200
rect 24044 24197 24072 24228
rect 24670 24216 24676 24268
rect 24728 24256 24734 24268
rect 25317 24259 25375 24265
rect 25317 24256 25329 24259
rect 24728 24228 25329 24256
rect 24728 24216 24734 24228
rect 25317 24225 25329 24228
rect 25363 24225 25375 24259
rect 25317 24219 25375 24225
rect 26326 24216 26332 24268
rect 26384 24256 26390 24268
rect 27433 24259 27491 24265
rect 27433 24256 27445 24259
rect 26384 24228 27445 24256
rect 26384 24216 26390 24228
rect 27433 24225 27445 24228
rect 27479 24225 27491 24259
rect 27433 24219 27491 24225
rect 23293 24191 23351 24197
rect 23293 24157 23305 24191
rect 23339 24188 23351 24191
rect 24029 24191 24087 24197
rect 23339 24160 23980 24188
rect 23339 24157 23351 24160
rect 23293 24151 23351 24157
rect 17052 24092 21036 24120
rect 21913 24123 21971 24129
rect 21913 24089 21925 24123
rect 21959 24089 21971 24123
rect 23753 24123 23811 24129
rect 23753 24120 23765 24123
rect 21913 24083 21971 24089
rect 22388 24092 23765 24120
rect 18230 24052 18236 24064
rect 18191 24024 18236 24052
rect 18230 24012 18236 24024
rect 18288 24012 18294 24064
rect 21928 24052 21956 24083
rect 22388 24064 22416 24092
rect 23753 24089 23765 24092
rect 23799 24120 23811 24123
rect 23842 24120 23848 24132
rect 23799 24092 23848 24120
rect 23799 24089 23811 24092
rect 23753 24083 23811 24089
rect 23842 24080 23848 24092
rect 23900 24080 23906 24132
rect 23952 24120 23980 24160
rect 24029 24157 24041 24191
rect 24075 24157 24087 24191
rect 24578 24188 24584 24200
rect 24539 24160 24584 24188
rect 24029 24151 24087 24157
rect 24578 24148 24584 24160
rect 24636 24148 24642 24200
rect 24762 24188 24768 24200
rect 24723 24160 24768 24188
rect 24762 24148 24768 24160
rect 24820 24148 24826 24200
rect 25406 24148 25412 24200
rect 25464 24188 25470 24200
rect 25573 24191 25631 24197
rect 25573 24188 25585 24191
rect 25464 24160 25585 24188
rect 25464 24148 25470 24160
rect 25573 24157 25585 24160
rect 25619 24157 25631 24191
rect 25573 24151 25631 24157
rect 27157 24191 27215 24197
rect 27157 24157 27169 24191
rect 27203 24188 27215 24191
rect 27614 24188 27620 24200
rect 27203 24160 27620 24188
rect 27203 24157 27215 24160
rect 27157 24151 27215 24157
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 28718 24188 28724 24200
rect 28679 24160 28724 24188
rect 28718 24148 28724 24160
rect 28776 24148 28782 24200
rect 28997 24191 29055 24197
rect 28997 24157 29009 24191
rect 29043 24188 29055 24191
rect 29270 24188 29276 24200
rect 29043 24160 29276 24188
rect 29043 24157 29055 24160
rect 28997 24151 29055 24157
rect 29270 24148 29276 24160
rect 29328 24188 29334 24200
rect 29932 24197 29960 24296
rect 31754 24256 31760 24268
rect 30760 24228 31760 24256
rect 30760 24197 30788 24228
rect 31754 24216 31760 24228
rect 31812 24216 31818 24268
rect 33428 24256 33456 24352
rect 33873 24259 33931 24265
rect 33873 24256 33885 24259
rect 33428 24228 33885 24256
rect 33873 24225 33885 24228
rect 33919 24225 33931 24259
rect 36170 24256 36176 24268
rect 36131 24228 36176 24256
rect 33873 24219 33931 24225
rect 36170 24216 36176 24228
rect 36228 24216 36234 24268
rect 29733 24191 29791 24197
rect 29733 24188 29745 24191
rect 29328 24160 29745 24188
rect 29328 24148 29334 24160
rect 29733 24157 29745 24160
rect 29779 24157 29791 24191
rect 29733 24151 29791 24157
rect 29917 24191 29975 24197
rect 29917 24157 29929 24191
rect 29963 24157 29975 24191
rect 29917 24151 29975 24157
rect 30653 24191 30711 24197
rect 30653 24157 30665 24191
rect 30699 24157 30711 24191
rect 30653 24151 30711 24157
rect 30745 24191 30803 24197
rect 30745 24157 30757 24191
rect 30791 24157 30803 24191
rect 30745 24151 30803 24157
rect 30929 24191 30987 24197
rect 30929 24157 30941 24191
rect 30975 24188 30987 24191
rect 31573 24191 31631 24197
rect 31573 24188 31585 24191
rect 30975 24160 31585 24188
rect 30975 24157 30987 24160
rect 30929 24151 30987 24157
rect 31573 24157 31585 24160
rect 31619 24157 31631 24191
rect 32030 24188 32036 24200
rect 31991 24160 32036 24188
rect 31573 24151 31631 24157
rect 24780 24120 24808 24148
rect 23952 24092 24808 24120
rect 30668 24120 30696 24151
rect 32030 24148 32036 24160
rect 32088 24148 32094 24200
rect 32122 24148 32128 24200
rect 32180 24188 32186 24200
rect 32289 24191 32347 24197
rect 32289 24188 32301 24191
rect 32180 24160 32301 24188
rect 32180 24148 32186 24160
rect 32289 24157 32301 24160
rect 32335 24157 32347 24191
rect 32289 24151 32347 24157
rect 34057 24191 34115 24197
rect 34057 24157 34069 24191
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34241 24191 34299 24197
rect 34241 24157 34253 24191
rect 34287 24188 34299 24191
rect 35069 24191 35127 24197
rect 35069 24188 35081 24191
rect 34287 24160 35081 24188
rect 34287 24157 34299 24160
rect 34241 24151 34299 24157
rect 35069 24157 35081 24160
rect 35115 24157 35127 24191
rect 35069 24151 35127 24157
rect 33870 24120 33876 24132
rect 30668 24092 33876 24120
rect 33870 24080 33876 24092
rect 33928 24080 33934 24132
rect 22370 24052 22376 24064
rect 21928 24024 22376 24052
rect 22370 24012 22376 24024
rect 22428 24012 22434 24064
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 23937 24055 23995 24061
rect 23937 24052 23949 24055
rect 22520 24024 23949 24052
rect 22520 24012 22526 24024
rect 23937 24021 23949 24024
rect 23983 24021 23995 24055
rect 31386 24052 31392 24064
rect 31347 24024 31392 24052
rect 23937 24015 23995 24021
rect 31386 24012 31392 24024
rect 31444 24012 31450 24064
rect 31754 24012 31760 24064
rect 31812 24052 31818 24064
rect 34072 24052 34100 24151
rect 36440 24123 36498 24129
rect 36440 24089 36452 24123
rect 36486 24120 36498 24123
rect 36630 24120 36636 24132
rect 36486 24092 36636 24120
rect 36486 24089 36498 24092
rect 36440 24083 36498 24089
rect 36630 24080 36636 24092
rect 36688 24080 36694 24132
rect 31812 24024 34100 24052
rect 31812 24012 31818 24024
rect 34790 24012 34796 24064
rect 34848 24052 34854 24064
rect 34885 24055 34943 24061
rect 34885 24052 34897 24055
rect 34848 24024 34897 24052
rect 34848 24012 34854 24024
rect 34885 24021 34897 24024
rect 34931 24021 34943 24055
rect 34885 24015 34943 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 17218 23808 17224 23860
rect 17276 23848 17282 23860
rect 17957 23851 18015 23857
rect 17957 23848 17969 23851
rect 17276 23820 17969 23848
rect 17276 23808 17282 23820
rect 17957 23817 17969 23820
rect 18003 23817 18015 23851
rect 17957 23811 18015 23817
rect 19429 23851 19487 23857
rect 19429 23817 19441 23851
rect 19475 23848 19487 23851
rect 19978 23848 19984 23860
rect 19475 23820 19984 23848
rect 19475 23817 19487 23820
rect 19429 23811 19487 23817
rect 19978 23808 19984 23820
rect 20036 23808 20042 23860
rect 21634 23808 21640 23860
rect 21692 23848 21698 23860
rect 22741 23851 22799 23857
rect 22741 23848 22753 23851
rect 21692 23820 22753 23848
rect 21692 23808 21698 23820
rect 22741 23817 22753 23820
rect 22787 23817 22799 23851
rect 22741 23811 22799 23817
rect 28718 23808 28724 23860
rect 28776 23848 28782 23860
rect 29089 23851 29147 23857
rect 29089 23848 29101 23851
rect 28776 23820 29101 23848
rect 28776 23808 28782 23820
rect 29089 23817 29101 23820
rect 29135 23817 29147 23851
rect 29089 23811 29147 23817
rect 29178 23808 29184 23860
rect 29236 23808 29242 23860
rect 32858 23808 32864 23860
rect 32916 23848 32922 23860
rect 36630 23848 36636 23860
rect 32916 23820 33088 23848
rect 36591 23820 36636 23848
rect 32916 23808 32922 23820
rect 17770 23740 17776 23792
rect 17828 23780 17834 23792
rect 17865 23783 17923 23789
rect 17865 23780 17877 23783
rect 17828 23752 17877 23780
rect 17828 23740 17834 23752
rect 17865 23749 17877 23752
rect 17911 23780 17923 23783
rect 23382 23780 23388 23792
rect 17911 23752 21404 23780
rect 23343 23752 23388 23780
rect 17911 23749 17923 23752
rect 17865 23743 17923 23749
rect 18230 23672 18236 23724
rect 18288 23712 18294 23724
rect 19245 23715 19303 23721
rect 19245 23712 19257 23715
rect 18288 23684 19257 23712
rect 18288 23672 18294 23684
rect 19245 23681 19257 23684
rect 19291 23681 19303 23715
rect 19426 23712 19432 23724
rect 19387 23684 19432 23712
rect 19245 23675 19303 23681
rect 19426 23672 19432 23684
rect 19484 23672 19490 23724
rect 21266 23712 21272 23724
rect 21227 23684 21272 23712
rect 21266 23672 21272 23684
rect 21324 23672 21330 23724
rect 21376 23712 21404 23752
rect 23382 23740 23388 23752
rect 23440 23740 23446 23792
rect 29196 23780 29224 23808
rect 29012 23752 29224 23780
rect 30460 23783 30518 23789
rect 22002 23712 22008 23724
rect 21376 23684 21772 23712
rect 21963 23684 22008 23712
rect 21744 23576 21772 23684
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 22186 23712 22192 23724
rect 22147 23684 22192 23712
rect 22186 23672 22192 23684
rect 22244 23672 22250 23724
rect 22370 23712 22376 23724
rect 22331 23684 22376 23712
rect 22370 23672 22376 23684
rect 22428 23672 22434 23724
rect 22554 23712 22560 23724
rect 22515 23684 22560 23712
rect 22554 23672 22560 23684
rect 22612 23672 22618 23724
rect 25958 23712 25964 23724
rect 25919 23684 25964 23712
rect 25958 23672 25964 23684
rect 26016 23672 26022 23724
rect 26053 23715 26111 23721
rect 26053 23681 26065 23715
rect 26099 23712 26111 23715
rect 26234 23712 26240 23724
rect 26099 23684 26240 23712
rect 26099 23681 26111 23684
rect 26053 23675 26111 23681
rect 26234 23672 26240 23684
rect 26292 23672 26298 23724
rect 26329 23715 26387 23721
rect 26329 23681 26341 23715
rect 26375 23712 26387 23715
rect 26970 23712 26976 23724
rect 26375 23684 26976 23712
rect 26375 23681 26387 23684
rect 26329 23675 26387 23681
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 29012 23721 29040 23752
rect 30460 23749 30472 23783
rect 30506 23780 30518 23783
rect 31386 23780 31392 23792
rect 30506 23752 31392 23780
rect 30506 23749 30518 23752
rect 30460 23743 30518 23749
rect 31386 23740 31392 23752
rect 31444 23740 31450 23792
rect 32950 23780 32956 23792
rect 32876 23752 32956 23780
rect 28997 23715 29055 23721
rect 28997 23681 29009 23715
rect 29043 23681 29055 23715
rect 28997 23675 29055 23681
rect 29181 23715 29239 23721
rect 29181 23681 29193 23715
rect 29227 23712 29239 23715
rect 29454 23712 29460 23724
rect 29227 23684 29460 23712
rect 29227 23681 29239 23684
rect 29181 23675 29239 23681
rect 29454 23672 29460 23684
rect 29512 23672 29518 23724
rect 32030 23712 32036 23724
rect 30208 23684 32036 23712
rect 21818 23604 21824 23656
rect 21876 23644 21882 23656
rect 22281 23647 22339 23653
rect 22281 23644 22293 23647
rect 21876 23616 22293 23644
rect 21876 23604 21882 23616
rect 22281 23613 22293 23616
rect 22327 23613 22339 23647
rect 25777 23647 25835 23653
rect 25777 23644 25789 23647
rect 22281 23607 22339 23613
rect 22572 23616 25789 23644
rect 22572 23576 22600 23616
rect 25777 23613 25789 23616
rect 25823 23613 25835 23647
rect 25777 23607 25835 23613
rect 29086 23604 29092 23656
rect 29144 23644 29150 23656
rect 30208 23653 30236 23684
rect 32030 23672 32036 23684
rect 32088 23672 32094 23724
rect 32876 23721 32904 23752
rect 32950 23740 32956 23752
rect 33008 23740 33014 23792
rect 33060 23721 33088 23820
rect 36630 23808 36636 23820
rect 36688 23808 36694 23860
rect 35526 23780 35532 23792
rect 35439 23752 35532 23780
rect 35526 23740 35532 23752
rect 35584 23780 35590 23792
rect 36170 23780 36176 23792
rect 35584 23752 36176 23780
rect 35584 23740 35590 23752
rect 36170 23740 36176 23752
rect 36228 23740 36234 23792
rect 32861 23715 32919 23721
rect 32861 23681 32873 23715
rect 32907 23681 32919 23715
rect 32861 23675 32919 23681
rect 33045 23715 33103 23721
rect 33045 23681 33057 23715
rect 33091 23681 33103 23715
rect 33778 23712 33784 23724
rect 33739 23684 33784 23712
rect 33045 23675 33103 23681
rect 33778 23672 33784 23684
rect 33836 23672 33842 23724
rect 36817 23715 36875 23721
rect 36817 23681 36829 23715
rect 36863 23712 36875 23715
rect 37274 23712 37280 23724
rect 36863 23684 37280 23712
rect 36863 23681 36875 23684
rect 36817 23675 36875 23681
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 37458 23712 37464 23724
rect 37419 23684 37464 23712
rect 37458 23672 37464 23684
rect 37516 23672 37522 23724
rect 37642 23712 37648 23724
rect 37603 23684 37648 23712
rect 37642 23672 37648 23684
rect 37700 23672 37706 23724
rect 30193 23647 30251 23653
rect 30193 23644 30205 23647
rect 29144 23616 30205 23644
rect 29144 23604 29150 23616
rect 30193 23613 30205 23616
rect 30239 23613 30251 23647
rect 30193 23607 30251 23613
rect 32769 23647 32827 23653
rect 32769 23613 32781 23647
rect 32815 23613 32827 23647
rect 32769 23607 32827 23613
rect 32953 23647 33011 23653
rect 32953 23613 32965 23647
rect 32999 23644 33011 23647
rect 33410 23644 33416 23656
rect 32999 23616 33416 23644
rect 32999 23613 33011 23616
rect 32953 23607 33011 23613
rect 21744 23548 22600 23576
rect 22646 23536 22652 23588
rect 22704 23576 22710 23588
rect 24673 23579 24731 23585
rect 24673 23576 24685 23579
rect 22704 23548 24685 23576
rect 22704 23536 22710 23548
rect 24673 23545 24685 23548
rect 24719 23545 24731 23579
rect 32784 23576 32812 23607
rect 33410 23604 33416 23616
rect 33468 23604 33474 23656
rect 34238 23576 34244 23588
rect 32784 23548 34244 23576
rect 24673 23539 24731 23545
rect 34238 23536 34244 23548
rect 34296 23536 34302 23588
rect 21361 23511 21419 23517
rect 21361 23477 21373 23511
rect 21407 23508 21419 23511
rect 21634 23508 21640 23520
rect 21407 23480 21640 23508
rect 21407 23477 21419 23480
rect 21361 23471 21419 23477
rect 21634 23468 21640 23480
rect 21692 23468 21698 23520
rect 26234 23508 26240 23520
rect 26195 23480 26240 23508
rect 26234 23468 26240 23480
rect 26292 23468 26298 23520
rect 31573 23511 31631 23517
rect 31573 23477 31585 23511
rect 31619 23508 31631 23511
rect 31938 23508 31944 23520
rect 31619 23480 31944 23508
rect 31619 23477 31631 23480
rect 31573 23471 31631 23477
rect 31938 23468 31944 23480
rect 31996 23468 32002 23520
rect 32582 23508 32588 23520
rect 32543 23480 32588 23508
rect 32582 23468 32588 23480
rect 32640 23468 32646 23520
rect 37550 23468 37556 23520
rect 37608 23508 37614 23520
rect 37829 23511 37887 23517
rect 37829 23508 37841 23511
rect 37608 23480 37841 23508
rect 37608 23468 37614 23480
rect 37829 23477 37841 23480
rect 37875 23477 37887 23511
rect 37829 23471 37887 23477
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 19426 23264 19432 23316
rect 19484 23304 19490 23316
rect 19613 23307 19671 23313
rect 19613 23304 19625 23307
rect 19484 23276 19625 23304
rect 19484 23264 19490 23276
rect 19613 23273 19625 23276
rect 19659 23304 19671 23307
rect 20438 23304 20444 23316
rect 19659 23276 20444 23304
rect 19659 23273 19671 23276
rect 19613 23267 19671 23273
rect 20438 23264 20444 23276
rect 20496 23264 20502 23316
rect 21361 23307 21419 23313
rect 21361 23273 21373 23307
rect 21407 23304 21419 23307
rect 22002 23304 22008 23316
rect 21407 23276 22008 23304
rect 21407 23273 21419 23276
rect 21361 23267 21419 23273
rect 22002 23264 22008 23276
rect 22060 23264 22066 23316
rect 23842 23264 23848 23316
rect 23900 23304 23906 23316
rect 24029 23307 24087 23313
rect 24029 23304 24041 23307
rect 23900 23276 24041 23304
rect 23900 23264 23906 23276
rect 24029 23273 24041 23276
rect 24075 23273 24087 23307
rect 25869 23307 25927 23313
rect 25869 23304 25881 23307
rect 24029 23267 24087 23273
rect 24136 23276 25881 23304
rect 20806 23168 20812 23180
rect 20767 23140 20812 23168
rect 20806 23128 20812 23140
rect 20864 23128 20870 23180
rect 22646 23168 22652 23180
rect 22607 23140 22652 23168
rect 22646 23128 22652 23140
rect 22704 23128 22710 23180
rect 17770 23100 17776 23112
rect 17731 23072 17776 23100
rect 17770 23060 17776 23072
rect 17828 23060 17834 23112
rect 17957 23103 18015 23109
rect 17957 23069 17969 23103
rect 18003 23100 18015 23103
rect 18003 23072 19288 23100
rect 18003 23069 18015 23072
rect 17957 23063 18015 23069
rect 17788 23032 17816 23060
rect 18632 23044 18660 23072
rect 18417 23035 18475 23041
rect 18417 23032 18429 23035
rect 17788 23004 18429 23032
rect 18417 23001 18429 23004
rect 18463 23001 18475 23035
rect 18417 22995 18475 23001
rect 18598 22992 18604 23044
rect 18656 23032 18662 23044
rect 19260 23032 19288 23072
rect 19334 23060 19340 23112
rect 19392 23100 19398 23112
rect 19429 23103 19487 23109
rect 19429 23100 19441 23103
rect 19392 23072 19441 23100
rect 19392 23060 19398 23072
rect 19429 23069 19441 23072
rect 19475 23100 19487 23103
rect 19978 23100 19984 23112
rect 19475 23072 19984 23100
rect 19475 23069 19487 23072
rect 19429 23063 19487 23069
rect 19978 23060 19984 23072
rect 20036 23060 20042 23112
rect 20714 23100 20720 23112
rect 20675 23072 20720 23100
rect 20714 23060 20720 23072
rect 20772 23060 20778 23112
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21266 23032 21272 23044
rect 18656 23004 18749 23032
rect 19260 23004 21272 23032
rect 18656 22992 18662 23004
rect 21266 22992 21272 23004
rect 21324 22992 21330 23044
rect 21560 23032 21588 23063
rect 21634 23060 21640 23112
rect 21692 23100 21698 23112
rect 21818 23100 21824 23112
rect 21692 23072 21737 23100
rect 21779 23072 21824 23100
rect 21692 23060 21698 23072
rect 21818 23060 21824 23072
rect 21876 23060 21882 23112
rect 21910 23060 21916 23112
rect 21968 23109 21974 23112
rect 21968 23103 21981 23109
rect 21969 23100 21981 23103
rect 21969 23072 22013 23100
rect 21969 23069 21981 23072
rect 21968 23063 21981 23069
rect 21968 23060 21974 23063
rect 22186 23032 22192 23044
rect 21560 23004 22192 23032
rect 22186 22992 22192 23004
rect 22244 22992 22250 23044
rect 22922 23041 22928 23044
rect 22916 23032 22928 23041
rect 22883 23004 22928 23032
rect 22916 22995 22928 23004
rect 22922 22992 22928 22995
rect 22980 22992 22986 23044
rect 17954 22964 17960 22976
rect 17915 22936 17960 22964
rect 17954 22924 17960 22936
rect 18012 22924 18018 22976
rect 18782 22964 18788 22976
rect 18743 22936 18788 22964
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 19334 22924 19340 22976
rect 19392 22964 19398 22976
rect 20254 22964 20260 22976
rect 19392 22936 20260 22964
rect 19392 22924 19398 22936
rect 20254 22924 20260 22936
rect 20312 22924 20318 22976
rect 21358 22924 21364 22976
rect 21416 22964 21422 22976
rect 24136 22964 24164 23276
rect 25869 23273 25881 23276
rect 25915 23273 25927 23307
rect 28997 23307 29055 23313
rect 28997 23304 29009 23307
rect 25869 23267 25927 23273
rect 26896 23276 29009 23304
rect 26896 23236 26924 23276
rect 28997 23273 29009 23276
rect 29043 23273 29055 23307
rect 31202 23304 31208 23316
rect 31163 23276 31208 23304
rect 28997 23267 29055 23273
rect 31202 23264 31208 23276
rect 31260 23304 31266 23316
rect 33778 23304 33784 23316
rect 31260 23276 33784 23304
rect 31260 23264 31266 23276
rect 33778 23264 33784 23276
rect 33836 23264 33842 23316
rect 34057 23307 34115 23313
rect 34057 23273 34069 23307
rect 34103 23273 34115 23307
rect 34238 23304 34244 23316
rect 34199 23276 34244 23304
rect 34057 23267 34115 23273
rect 32306 23236 32312 23248
rect 25148 23208 26924 23236
rect 32267 23208 32312 23236
rect 25148 23109 25176 23208
rect 25317 23171 25375 23177
rect 25317 23137 25329 23171
rect 25363 23168 25375 23171
rect 26234 23168 26240 23180
rect 25363 23140 26240 23168
rect 25363 23137 25375 23140
rect 25317 23131 25375 23137
rect 26068 23109 26096 23140
rect 26234 23128 26240 23140
rect 26292 23128 26298 23180
rect 26326 23128 26332 23180
rect 26384 23168 26390 23180
rect 26384 23140 26429 23168
rect 26384 23128 26390 23140
rect 25041 23103 25099 23109
rect 25041 23069 25053 23103
rect 25087 23069 25099 23103
rect 25041 23063 25099 23069
rect 25133 23103 25191 23109
rect 25133 23069 25145 23103
rect 25179 23069 25191 23103
rect 25133 23063 25191 23069
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23069 26111 23103
rect 26053 23063 26111 23069
rect 26145 23103 26203 23109
rect 26145 23069 26157 23103
rect 26191 23069 26203 23103
rect 26145 23063 26203 23069
rect 26421 23103 26479 23109
rect 26421 23069 26433 23103
rect 26467 23100 26479 23103
rect 26786 23100 26792 23112
rect 26467 23072 26792 23100
rect 26467 23069 26479 23072
rect 26421 23063 26479 23069
rect 25056 23032 25084 23063
rect 25056 23004 25728 23032
rect 25700 22976 25728 23004
rect 25958 22992 25964 23044
rect 26016 23032 26022 23044
rect 26160 23032 26188 23063
rect 26786 23060 26792 23072
rect 26844 23060 26850 23112
rect 26896 23109 26924 23208
rect 32306 23196 32312 23208
rect 32364 23196 32370 23248
rect 32769 23239 32827 23245
rect 32769 23205 32781 23239
rect 32815 23236 32827 23239
rect 32858 23236 32864 23248
rect 32815 23208 32864 23236
rect 32815 23205 32827 23208
rect 32769 23199 32827 23205
rect 32858 23196 32864 23208
rect 32916 23196 32922 23248
rect 31938 23168 31944 23180
rect 31851 23140 31944 23168
rect 31938 23128 31944 23140
rect 31996 23168 32002 23180
rect 34072 23168 34100 23267
rect 34238 23264 34244 23276
rect 34296 23264 34302 23316
rect 38286 23304 38292 23316
rect 38247 23276 38292 23304
rect 38286 23264 38292 23276
rect 38344 23264 38350 23316
rect 31996 23140 34100 23168
rect 31996 23128 32002 23140
rect 36170 23128 36176 23180
rect 36228 23168 36234 23180
rect 36909 23171 36967 23177
rect 36909 23168 36921 23171
rect 36228 23140 36921 23168
rect 36228 23128 36234 23140
rect 36909 23137 36921 23140
rect 36955 23137 36967 23171
rect 36909 23131 36967 23137
rect 26881 23103 26939 23109
rect 26881 23069 26893 23103
rect 26927 23069 26939 23103
rect 26881 23063 26939 23069
rect 27065 23103 27123 23109
rect 27065 23069 27077 23103
rect 27111 23069 27123 23103
rect 27065 23063 27123 23069
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 28994 23100 29000 23112
rect 27663 23072 29000 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 26973 23035 27031 23041
rect 26973 23032 26985 23035
rect 26016 23004 26985 23032
rect 26016 22992 26022 23004
rect 26973 23001 26985 23004
rect 27019 23001 27031 23035
rect 26973 22995 27031 23001
rect 21416 22936 24164 22964
rect 21416 22924 21422 22936
rect 25682 22924 25688 22976
rect 25740 22964 25746 22976
rect 27080 22964 27108 23063
rect 28994 23060 29000 23072
rect 29052 23060 29058 23112
rect 31754 23060 31760 23112
rect 31812 23100 31818 23112
rect 32125 23103 32183 23109
rect 32125 23100 32137 23103
rect 31812 23072 32137 23100
rect 31812 23060 31818 23072
rect 32125 23069 32137 23072
rect 32171 23069 32183 23103
rect 33042 23100 33048 23112
rect 33003 23072 33048 23100
rect 32125 23063 32183 23069
rect 33042 23060 33048 23072
rect 33100 23060 33106 23112
rect 33137 23103 33195 23109
rect 33137 23078 33149 23103
rect 33183 23078 33195 23103
rect 33234 23103 33292 23109
rect 27884 23035 27942 23041
rect 27884 23001 27896 23035
rect 27930 23032 27942 23035
rect 29086 23032 29092 23044
rect 27930 23004 29092 23032
rect 27930 23001 27942 23004
rect 27884 22995 27942 23001
rect 29086 22992 29092 23004
rect 29144 22992 29150 23044
rect 29733 23035 29791 23041
rect 29733 23001 29745 23035
rect 29779 23032 29791 23035
rect 29779 23004 33088 23032
rect 33134 23026 33140 23078
rect 33192 23026 33198 23078
rect 33234 23069 33246 23103
rect 33280 23100 33292 23103
rect 33413 23103 33471 23109
rect 33280 23072 33364 23100
rect 33280 23069 33292 23072
rect 33234 23063 33292 23069
rect 33336 23032 33364 23072
rect 33413 23069 33425 23103
rect 33459 23100 33471 23103
rect 33502 23100 33508 23112
rect 33459 23072 33508 23100
rect 33459 23069 33471 23072
rect 33413 23063 33471 23069
rect 33502 23060 33508 23072
rect 33560 23060 33566 23112
rect 34882 23100 34888 23112
rect 34795 23072 34888 23100
rect 34882 23060 34888 23072
rect 34940 23100 34946 23112
rect 35526 23100 35532 23112
rect 34940 23072 35532 23100
rect 34940 23060 34946 23072
rect 35526 23060 35532 23072
rect 35584 23060 35590 23112
rect 33686 23032 33692 23044
rect 33336 23004 33692 23032
rect 29779 23001 29791 23004
rect 29733 22995 29791 23001
rect 25740 22936 27108 22964
rect 33060 22964 33088 23004
rect 33686 22992 33692 23004
rect 33744 22992 33750 23044
rect 33870 23032 33876 23044
rect 33831 23004 33876 23032
rect 33870 22992 33876 23004
rect 33928 22992 33934 23044
rect 34514 23032 34520 23044
rect 33980 23004 34520 23032
rect 33980 22964 34008 23004
rect 34514 22992 34520 23004
rect 34572 22992 34578 23044
rect 34790 22992 34796 23044
rect 34848 23032 34854 23044
rect 35130 23035 35188 23041
rect 35130 23032 35142 23035
rect 34848 23004 35142 23032
rect 34848 22992 34854 23004
rect 35130 23001 35142 23004
rect 35176 23001 35188 23035
rect 35130 22995 35188 23001
rect 37176 23035 37234 23041
rect 37176 23001 37188 23035
rect 37222 23032 37234 23035
rect 37366 23032 37372 23044
rect 37222 23004 37372 23032
rect 37222 23001 37234 23004
rect 37176 22995 37234 23001
rect 37366 22992 37372 23004
rect 37424 22992 37430 23044
rect 33060 22936 34008 22964
rect 34083 22967 34141 22973
rect 25740 22924 25746 22936
rect 34083 22933 34095 22967
rect 34129 22964 34141 22967
rect 35526 22964 35532 22976
rect 34129 22936 35532 22964
rect 34129 22933 34141 22936
rect 34083 22927 34141 22933
rect 35526 22924 35532 22936
rect 35584 22924 35590 22976
rect 35802 22924 35808 22976
rect 35860 22964 35866 22976
rect 36265 22967 36323 22973
rect 36265 22964 36277 22967
rect 35860 22936 36277 22964
rect 35860 22924 35866 22936
rect 36265 22933 36277 22936
rect 36311 22933 36323 22967
rect 36265 22927 36323 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 17862 22760 17868 22772
rect 17823 22732 17868 22760
rect 17862 22720 17868 22732
rect 17920 22720 17926 22772
rect 17957 22763 18015 22769
rect 17957 22729 17969 22763
rect 18003 22760 18015 22763
rect 18046 22760 18052 22772
rect 18003 22732 18052 22760
rect 18003 22729 18015 22732
rect 17957 22723 18015 22729
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 18782 22760 18788 22772
rect 18340 22732 18788 22760
rect 17589 22627 17647 22633
rect 17589 22593 17601 22627
rect 17635 22624 17647 22627
rect 17954 22624 17960 22636
rect 17635 22596 17960 22624
rect 17635 22593 17647 22596
rect 17589 22587 17647 22593
rect 17954 22584 17960 22596
rect 18012 22584 18018 22636
rect 18049 22627 18107 22633
rect 18049 22593 18061 22627
rect 18095 22624 18107 22627
rect 18138 22624 18144 22636
rect 18095 22596 18144 22624
rect 18095 22593 18107 22596
rect 18049 22587 18107 22593
rect 18138 22584 18144 22596
rect 18196 22624 18202 22636
rect 18340 22624 18368 22732
rect 18782 22720 18788 22732
rect 18840 22720 18846 22772
rect 19426 22760 19432 22772
rect 18892 22732 19432 22760
rect 18892 22639 18920 22732
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 20993 22763 21051 22769
rect 20993 22729 21005 22763
rect 21039 22760 21051 22763
rect 21266 22760 21272 22772
rect 21039 22732 21272 22760
rect 21039 22729 21051 22732
rect 20993 22723 21051 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 21818 22720 21824 22772
rect 21876 22760 21882 22772
rect 21876 22732 22816 22760
rect 21876 22720 21882 22732
rect 19858 22695 19916 22701
rect 19858 22692 19870 22695
rect 19306 22664 19870 22692
rect 18196 22596 18368 22624
rect 18196 22584 18202 22596
rect 18598 22584 18604 22636
rect 18656 22628 18662 22636
rect 18874 22633 18932 22639
rect 18785 22628 18843 22633
rect 18656 22627 18843 22628
rect 18656 22600 18797 22627
rect 18656 22584 18662 22600
rect 18785 22593 18797 22600
rect 18831 22593 18843 22627
rect 18874 22599 18886 22633
rect 18920 22599 18932 22633
rect 18874 22593 18932 22599
rect 18969 22630 19027 22636
rect 18969 22596 18981 22630
rect 19015 22596 19027 22630
rect 19150 22624 19156 22636
rect 19111 22596 19156 22624
rect 18785 22587 18843 22593
rect 18969 22590 19027 22596
rect 18984 22556 19012 22590
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19058 22556 19064 22568
rect 18984 22528 19064 22556
rect 19058 22516 19064 22528
rect 19116 22516 19122 22568
rect 18509 22491 18567 22497
rect 18509 22457 18521 22491
rect 18555 22488 18567 22491
rect 19306 22488 19334 22664
rect 19858 22661 19870 22664
rect 19904 22661 19916 22695
rect 19858 22655 19916 22661
rect 22370 22652 22376 22704
rect 22428 22692 22434 22704
rect 22788 22701 22816 22732
rect 22922 22720 22928 22772
rect 22980 22760 22986 22772
rect 23385 22763 23443 22769
rect 23385 22760 23397 22763
rect 22980 22732 23397 22760
rect 22980 22720 22986 22732
rect 23385 22729 23397 22732
rect 23431 22729 23443 22763
rect 25682 22760 25688 22772
rect 25643 22732 25688 22760
rect 23385 22723 23443 22729
rect 25682 22720 25688 22732
rect 25740 22720 25746 22772
rect 26326 22720 26332 22772
rect 26384 22760 26390 22772
rect 26605 22763 26663 22769
rect 26605 22760 26617 22763
rect 26384 22732 26617 22760
rect 26384 22720 26390 22732
rect 26605 22729 26617 22732
rect 26651 22729 26663 22763
rect 30558 22760 30564 22772
rect 30519 22732 30564 22760
rect 26605 22723 26663 22729
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 33686 22760 33692 22772
rect 33647 22732 33692 22760
rect 33686 22720 33692 22732
rect 33744 22760 33750 22772
rect 33962 22760 33968 22772
rect 33744 22732 33968 22760
rect 33744 22720 33750 22732
rect 33962 22720 33968 22732
rect 34020 22720 34026 22772
rect 34241 22763 34299 22769
rect 34241 22729 34253 22763
rect 34287 22729 34299 22763
rect 34241 22723 34299 22729
rect 22557 22695 22615 22701
rect 22557 22692 22569 22695
rect 22428 22664 22569 22692
rect 22428 22652 22434 22664
rect 22557 22661 22569 22664
rect 22603 22661 22615 22695
rect 22557 22655 22615 22661
rect 22773 22695 22831 22701
rect 22773 22661 22785 22695
rect 22819 22692 22831 22695
rect 23566 22692 23572 22704
rect 22819 22664 23572 22692
rect 22819 22661 22831 22664
rect 22773 22655 22831 22661
rect 23566 22652 23572 22664
rect 23624 22652 23630 22704
rect 23661 22695 23719 22701
rect 23661 22661 23673 22695
rect 23707 22692 23719 22695
rect 24026 22692 24032 22704
rect 23707 22664 24032 22692
rect 23707 22661 23719 22664
rect 23661 22655 23719 22661
rect 24026 22652 24032 22664
rect 24084 22692 24090 22704
rect 24394 22692 24400 22704
rect 24084 22664 24400 22692
rect 24084 22652 24090 22664
rect 24394 22652 24400 22664
rect 24452 22652 24458 22704
rect 31110 22692 31116 22704
rect 29748 22664 31116 22692
rect 23106 22584 23112 22636
rect 23164 22624 23170 22636
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23164 22596 23397 22624
rect 23164 22584 23170 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 23477 22627 23535 22633
rect 23477 22593 23489 22627
rect 23523 22624 23535 22627
rect 23750 22624 23756 22636
rect 23523 22596 23756 22624
rect 23523 22593 23535 22596
rect 23477 22587 23535 22593
rect 23750 22584 23756 22596
rect 23808 22584 23814 22636
rect 24578 22633 24584 22636
rect 24572 22587 24584 22633
rect 24636 22624 24642 22636
rect 27982 22633 27988 22636
rect 24636 22596 24672 22624
rect 24578 22584 24584 22587
rect 24636 22584 24642 22596
rect 27976 22587 27988 22633
rect 28040 22624 28046 22636
rect 29748 22633 29776 22664
rect 31110 22652 31116 22664
rect 31168 22652 31174 22704
rect 32582 22701 32588 22704
rect 32576 22692 32588 22701
rect 32543 22664 32588 22692
rect 32576 22655 32588 22664
rect 32582 22652 32588 22655
rect 32640 22652 32646 22704
rect 34256 22692 34284 22723
rect 37274 22720 37280 22772
rect 37332 22760 37338 22772
rect 37829 22763 37887 22769
rect 37829 22760 37841 22763
rect 37332 22732 37841 22760
rect 37332 22720 37338 22732
rect 37829 22729 37841 22732
rect 37875 22729 37887 22763
rect 37829 22723 37887 22729
rect 35130 22695 35188 22701
rect 35130 22692 35142 22695
rect 34256 22664 35142 22692
rect 35130 22661 35142 22664
rect 35176 22661 35188 22695
rect 38286 22692 38292 22704
rect 35130 22655 35188 22661
rect 37568 22664 38292 22692
rect 29733 22627 29791 22633
rect 28040 22596 28076 22624
rect 27982 22584 27988 22587
rect 28040 22584 28046 22596
rect 29733 22593 29745 22627
rect 29779 22593 29791 22627
rect 30282 22624 30288 22636
rect 30243 22596 30288 22624
rect 29733 22587 29791 22593
rect 30282 22584 30288 22596
rect 30340 22584 30346 22636
rect 31297 22627 31355 22633
rect 31297 22593 31309 22627
rect 31343 22624 31355 22627
rect 31343 22596 31984 22624
rect 31343 22593 31355 22596
rect 31297 22587 31355 22593
rect 19426 22516 19432 22568
rect 19484 22556 19490 22568
rect 19613 22559 19671 22565
rect 19613 22556 19625 22559
rect 19484 22528 19625 22556
rect 19484 22516 19490 22528
rect 19613 22525 19625 22528
rect 19659 22525 19671 22559
rect 24302 22556 24308 22568
rect 24263 22528 24308 22556
rect 19613 22519 19671 22525
rect 24302 22516 24308 22528
rect 24360 22516 24366 22568
rect 25774 22516 25780 22568
rect 25832 22556 25838 22568
rect 26145 22559 26203 22565
rect 26145 22556 26157 22559
rect 25832 22528 26157 22556
rect 25832 22516 25838 22528
rect 26145 22525 26157 22528
rect 26191 22525 26203 22559
rect 26510 22556 26516 22568
rect 26423 22528 26516 22556
rect 26145 22519 26203 22525
rect 18555 22460 19334 22488
rect 22925 22491 22983 22497
rect 18555 22457 18567 22460
rect 18509 22451 18567 22457
rect 22925 22457 22937 22491
rect 22971 22488 22983 22491
rect 23106 22488 23112 22500
rect 22971 22460 23112 22488
rect 22971 22457 22983 22460
rect 22925 22451 22983 22457
rect 23106 22448 23112 22460
rect 23164 22448 23170 22500
rect 26436 22497 26464 22528
rect 26510 22516 26516 22528
rect 26568 22556 26574 22568
rect 27706 22556 27712 22568
rect 26568 22528 27292 22556
rect 27667 22528 27712 22556
rect 26568 22516 26574 22528
rect 26421 22491 26479 22497
rect 26421 22457 26433 22491
rect 26467 22457 26479 22491
rect 26421 22451 26479 22457
rect 19978 22380 19984 22432
rect 20036 22420 20042 22432
rect 21358 22420 21364 22432
rect 20036 22392 21364 22420
rect 20036 22380 20042 22392
rect 21358 22380 21364 22392
rect 21416 22380 21422 22432
rect 22186 22380 22192 22432
rect 22244 22420 22250 22432
rect 22554 22420 22560 22432
rect 22244 22392 22560 22420
rect 22244 22380 22250 22392
rect 22554 22380 22560 22392
rect 22612 22420 22618 22432
rect 22741 22423 22799 22429
rect 22741 22420 22753 22423
rect 22612 22392 22753 22420
rect 22612 22380 22618 22392
rect 22741 22389 22753 22392
rect 22787 22389 22799 22423
rect 27264 22420 27292 22528
rect 27706 22516 27712 22528
rect 27764 22516 27770 22568
rect 31113 22559 31171 22565
rect 31113 22556 31125 22559
rect 29104 22528 31125 22556
rect 29104 22497 29132 22528
rect 31113 22525 31125 22528
rect 31159 22525 31171 22559
rect 31113 22519 31171 22525
rect 29089 22491 29147 22497
rect 29089 22457 29101 22491
rect 29135 22457 29147 22491
rect 29089 22451 29147 22457
rect 29549 22491 29607 22497
rect 29549 22457 29561 22491
rect 29595 22488 29607 22491
rect 30558 22488 30564 22500
rect 29595 22460 30564 22488
rect 29595 22457 29607 22460
rect 29549 22451 29607 22457
rect 29104 22420 29132 22451
rect 30558 22448 30564 22460
rect 30616 22448 30622 22500
rect 31478 22420 31484 22432
rect 27264 22392 29132 22420
rect 31439 22392 31484 22420
rect 22741 22383 22799 22389
rect 31478 22380 31484 22392
rect 31536 22380 31542 22432
rect 31956 22420 31984 22596
rect 32030 22584 32036 22636
rect 32088 22624 32094 22636
rect 32309 22627 32367 22633
rect 32309 22624 32321 22627
rect 32088 22596 32321 22624
rect 32088 22584 32094 22596
rect 32309 22593 32321 22596
rect 32355 22593 32367 22627
rect 32309 22587 32367 22593
rect 33134 22584 33140 22636
rect 33192 22624 33198 22636
rect 34422 22624 34428 22636
rect 33192 22596 34284 22624
rect 34383 22596 34428 22624
rect 33192 22584 33198 22596
rect 33410 22420 33416 22432
rect 31956 22392 33416 22420
rect 33410 22380 33416 22392
rect 33468 22380 33474 22432
rect 34256 22420 34284 22596
rect 34422 22584 34428 22596
rect 34480 22584 34486 22636
rect 34882 22624 34888 22636
rect 34843 22596 34888 22624
rect 34882 22584 34888 22596
rect 34940 22584 34946 22636
rect 37568 22633 37596 22664
rect 38286 22652 38292 22664
rect 38344 22652 38350 22704
rect 37553 22627 37611 22633
rect 37553 22593 37565 22627
rect 37599 22593 37611 22627
rect 37553 22587 37611 22593
rect 37642 22584 37648 22636
rect 37700 22624 37706 22636
rect 37700 22596 37745 22624
rect 37700 22584 37706 22596
rect 35618 22420 35624 22432
rect 34256 22392 35624 22420
rect 35618 22380 35624 22392
rect 35676 22380 35682 22432
rect 36262 22420 36268 22432
rect 36223 22392 36268 22420
rect 36262 22380 36268 22392
rect 36320 22380 36326 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 18601 22219 18659 22225
rect 18601 22185 18613 22219
rect 18647 22216 18659 22219
rect 18782 22216 18788 22228
rect 18647 22188 18788 22216
rect 18647 22185 18659 22188
rect 18601 22179 18659 22185
rect 18782 22176 18788 22188
rect 18840 22176 18846 22228
rect 20438 22216 20444 22228
rect 20399 22188 20444 22216
rect 20438 22176 20444 22188
rect 20496 22176 20502 22228
rect 22465 22219 22523 22225
rect 22465 22185 22477 22219
rect 22511 22216 22523 22219
rect 22511 22188 23336 22216
rect 22511 22185 22523 22188
rect 22465 22179 22523 22185
rect 20993 22151 21051 22157
rect 20993 22117 21005 22151
rect 21039 22148 21051 22151
rect 23017 22151 23075 22157
rect 21039 22120 21073 22148
rect 21039 22117 21051 22120
rect 20993 22111 21051 22117
rect 23017 22117 23029 22151
rect 23063 22148 23075 22151
rect 23063 22120 23097 22148
rect 23063 22117 23075 22120
rect 23017 22111 23075 22117
rect 17753 22083 17811 22089
rect 17753 22049 17765 22083
rect 17799 22080 17811 22083
rect 17862 22080 17868 22092
rect 17799 22052 17868 22080
rect 17799 22049 17811 22052
rect 17753 22043 17811 22049
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 21008 22080 21036 22111
rect 23032 22080 23060 22111
rect 20272 22052 21036 22080
rect 22296 22052 23060 22080
rect 17954 22012 17960 22024
rect 17867 21984 17960 22012
rect 17954 21972 17960 21984
rect 18012 22012 18018 22024
rect 20272 22021 20300 22052
rect 20257 22015 20315 22021
rect 18012 21984 18552 22012
rect 18012 21972 18018 21984
rect 17681 21947 17739 21953
rect 17681 21913 17693 21947
rect 17727 21944 17739 21947
rect 17865 21947 17923 21953
rect 17727 21916 17816 21944
rect 17727 21913 17739 21916
rect 17681 21907 17739 21913
rect 17788 21876 17816 21916
rect 17865 21913 17877 21947
rect 17911 21944 17923 21947
rect 18138 21944 18144 21956
rect 17911 21916 18144 21944
rect 17911 21913 17923 21916
rect 17865 21907 17923 21913
rect 18138 21904 18144 21916
rect 18196 21904 18202 21956
rect 18417 21947 18475 21953
rect 18417 21913 18429 21947
rect 18463 21913 18475 21947
rect 18524 21944 18552 21984
rect 20257 21981 20269 22015
rect 20303 21981 20315 22015
rect 20257 21975 20315 21981
rect 20533 22015 20591 22021
rect 20533 21981 20545 22015
rect 20579 22012 20591 22015
rect 20714 22012 20720 22024
rect 20579 21984 20720 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 18617 21947 18675 21953
rect 18617 21944 18629 21947
rect 18524 21916 18629 21944
rect 18417 21907 18475 21913
rect 18617 21913 18629 21916
rect 18663 21913 18675 21947
rect 20548 21944 20576 21975
rect 20714 21972 20720 21984
rect 20772 22012 20778 22024
rect 21174 22012 21180 22024
rect 20772 21984 21180 22012
rect 20772 21972 20778 21984
rect 21174 21972 21180 21984
rect 21232 21972 21238 22024
rect 21269 22015 21327 22021
rect 21269 21981 21281 22015
rect 21315 22012 21327 22015
rect 21358 22012 21364 22024
rect 21315 21984 21364 22012
rect 21315 21981 21327 21984
rect 21269 21975 21327 21981
rect 21358 21972 21364 21984
rect 21416 21972 21422 22024
rect 22296 22021 22324 22052
rect 22281 22015 22339 22021
rect 22281 21981 22293 22015
rect 22327 21981 22339 22015
rect 22554 22012 22560 22024
rect 22467 21984 22560 22012
rect 22281 21975 22339 21981
rect 22554 21972 22560 21984
rect 22612 22012 22618 22024
rect 23106 22012 23112 22024
rect 22612 21984 23112 22012
rect 22612 21972 22618 21984
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23308 22021 23336 22188
rect 24578 22176 24584 22228
rect 24636 22216 24642 22228
rect 24765 22219 24823 22225
rect 24765 22216 24777 22219
rect 24636 22188 24777 22216
rect 24636 22176 24642 22188
rect 24765 22185 24777 22188
rect 24811 22185 24823 22219
rect 28997 22219 29055 22225
rect 24765 22179 24823 22185
rect 26896 22188 27568 22216
rect 26896 22157 26924 22188
rect 26881 22151 26939 22157
rect 26881 22148 26893 22151
rect 26791 22120 26893 22148
rect 26881 22117 26893 22120
rect 26927 22117 26939 22151
rect 26881 22111 26939 22117
rect 26053 22083 26111 22089
rect 26053 22080 26065 22083
rect 24964 22052 26065 22080
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 22012 23351 22015
rect 23566 22012 23572 22024
rect 23339 21984 23572 22012
rect 23339 21981 23351 21984
rect 23293 21975 23351 21981
rect 23566 21972 23572 21984
rect 23624 21972 23630 22024
rect 24964 22021 24992 22052
rect 26053 22049 26065 22052
rect 26099 22049 26111 22083
rect 26510 22080 26516 22092
rect 26471 22052 26516 22080
rect 26053 22043 26111 22049
rect 26510 22040 26516 22052
rect 26568 22040 26574 22092
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 25774 22012 25780 22024
rect 25687 21984 25780 22012
rect 24949 21975 25007 21981
rect 25774 21972 25780 21984
rect 25832 21972 25838 22024
rect 25869 22015 25927 22021
rect 25869 21981 25881 22015
rect 25915 22012 25927 22015
rect 26786 22012 26792 22024
rect 25915 21984 26792 22012
rect 25915 21981 25927 21984
rect 25869 21975 25927 21981
rect 26786 21972 26792 21984
rect 26844 21972 26850 22024
rect 18617 21907 18675 21913
rect 18708 21916 20576 21944
rect 18046 21876 18052 21888
rect 17788 21848 18052 21876
rect 18046 21836 18052 21848
rect 18104 21876 18110 21888
rect 18432 21876 18460 21907
rect 18708 21876 18736 21916
rect 20898 21904 20904 21956
rect 20956 21944 20962 21956
rect 20993 21947 21051 21953
rect 20993 21944 21005 21947
rect 20956 21916 21005 21944
rect 20956 21904 20962 21916
rect 20993 21913 21005 21916
rect 21039 21944 21051 21947
rect 23017 21947 23075 21953
rect 23017 21944 23029 21947
rect 21039 21916 23029 21944
rect 21039 21913 21051 21916
rect 20993 21907 21051 21913
rect 23017 21913 23029 21916
rect 23063 21944 23075 21947
rect 25222 21944 25228 21956
rect 23063 21916 25228 21944
rect 23063 21913 23075 21916
rect 23017 21907 23075 21913
rect 25222 21904 25228 21916
rect 25280 21904 25286 21956
rect 25792 21944 25820 21972
rect 26896 21944 26924 22111
rect 26970 22108 26976 22160
rect 27028 22148 27034 22160
rect 27028 22120 27073 22148
rect 27028 22108 27034 22120
rect 25792 21916 26924 21944
rect 18104 21848 18736 21876
rect 18785 21879 18843 21885
rect 18104 21836 18110 21848
rect 18785 21845 18797 21879
rect 18831 21876 18843 21879
rect 18874 21876 18880 21888
rect 18831 21848 18880 21876
rect 18831 21845 18843 21848
rect 18785 21839 18843 21845
rect 18874 21836 18880 21848
rect 18932 21836 18938 21888
rect 20070 21876 20076 21888
rect 20031 21848 20076 21876
rect 20070 21836 20076 21848
rect 20128 21836 20134 21888
rect 22094 21836 22100 21888
rect 22152 21876 22158 21888
rect 23198 21876 23204 21888
rect 22152 21848 22197 21876
rect 23159 21848 23204 21876
rect 22152 21836 22158 21848
rect 23198 21836 23204 21848
rect 23256 21836 23262 21888
rect 27540 21876 27568 22188
rect 28997 22185 29009 22219
rect 29043 22216 29055 22219
rect 29086 22216 29092 22228
rect 29043 22188 29092 22216
rect 29043 22185 29055 22188
rect 28997 22179 29055 22185
rect 29086 22176 29092 22188
rect 29144 22176 29150 22228
rect 31754 22176 31760 22228
rect 31812 22216 31818 22228
rect 33321 22219 33379 22225
rect 33321 22216 33333 22219
rect 31812 22188 33333 22216
rect 31812 22176 31818 22188
rect 33321 22185 33333 22188
rect 33367 22185 33379 22219
rect 33321 22179 33379 22185
rect 34333 22219 34391 22225
rect 34333 22185 34345 22219
rect 34379 22216 34391 22219
rect 34422 22216 34428 22228
rect 34379 22188 34428 22216
rect 34379 22185 34391 22188
rect 34333 22179 34391 22185
rect 28353 22151 28411 22157
rect 28353 22117 28365 22151
rect 28399 22148 28411 22151
rect 28399 22120 28856 22148
rect 28399 22117 28411 22120
rect 28353 22111 28411 22117
rect 28534 22012 28540 22024
rect 28495 21984 28540 22012
rect 28534 21972 28540 21984
rect 28592 21972 28598 22024
rect 28828 22012 28856 22120
rect 32401 22083 32459 22089
rect 32401 22049 32413 22083
rect 32447 22080 32459 22083
rect 33134 22080 33140 22092
rect 32447 22052 33140 22080
rect 32447 22049 32459 22052
rect 32401 22043 32459 22049
rect 33134 22040 33140 22052
rect 33192 22040 33198 22092
rect 33336 22080 33364 22179
rect 34422 22176 34428 22188
rect 34480 22176 34486 22228
rect 35158 22176 35164 22228
rect 35216 22216 35222 22228
rect 35802 22216 35808 22228
rect 35216 22188 35808 22216
rect 35216 22176 35222 22188
rect 35802 22176 35808 22188
rect 35860 22216 35866 22228
rect 35989 22219 36047 22225
rect 35989 22216 36001 22219
rect 35860 22188 36001 22216
rect 35860 22176 35866 22188
rect 35989 22185 36001 22188
rect 36035 22185 36047 22219
rect 37366 22216 37372 22228
rect 37327 22188 37372 22216
rect 35989 22179 36047 22185
rect 37366 22176 37372 22188
rect 37424 22176 37430 22228
rect 35386 22120 35664 22148
rect 33336 22052 34192 22080
rect 34164 22024 34192 22052
rect 34698 22040 34704 22092
rect 34756 22080 34762 22092
rect 34977 22083 35035 22089
rect 34977 22080 34989 22083
rect 34756 22052 34989 22080
rect 34756 22040 34762 22052
rect 34977 22049 34989 22052
rect 35023 22080 35035 22083
rect 35386 22080 35414 22120
rect 35526 22080 35532 22092
rect 35023 22052 35414 22080
rect 35487 22052 35532 22080
rect 35023 22049 35035 22052
rect 34977 22043 35035 22049
rect 35526 22040 35532 22052
rect 35584 22040 35590 22092
rect 35636 22080 35664 22120
rect 36170 22080 36176 22092
rect 35636 22052 36032 22080
rect 36131 22052 36176 22080
rect 28994 22012 29000 22024
rect 28828 21984 29000 22012
rect 28994 21972 29000 21984
rect 29052 21972 29058 22024
rect 29181 22015 29239 22021
rect 29181 21981 29193 22015
rect 29227 21981 29239 22015
rect 30006 22012 30012 22024
rect 29967 21984 30012 22012
rect 29181 21975 29239 21981
rect 29196 21944 29224 21975
rect 30006 21972 30012 21984
rect 30064 21972 30070 22024
rect 31478 22012 31484 22024
rect 30208 21984 31484 22012
rect 30208 21944 30236 21984
rect 31478 21972 31484 21984
rect 31536 21972 31542 22024
rect 32309 22015 32367 22021
rect 32309 21981 32321 22015
rect 32355 21981 32367 22015
rect 32490 22012 32496 22024
rect 32451 21984 32496 22012
rect 32309 21975 32367 21981
rect 29196 21916 30236 21944
rect 30276 21947 30334 21953
rect 30276 21913 30288 21947
rect 30322 21944 30334 21947
rect 32324 21944 32352 21975
rect 32490 21972 32496 21984
rect 32548 21972 32554 22024
rect 32582 21972 32588 22024
rect 32640 22012 32646 22024
rect 33594 22012 33600 22024
rect 32640 21984 32685 22012
rect 33152 21984 33600 22012
rect 32640 21972 32646 21984
rect 33152 21944 33180 21984
rect 33594 21972 33600 21984
rect 33652 21972 33658 22024
rect 34057 22015 34115 22021
rect 34057 21981 34069 22015
rect 34103 21981 34115 22015
rect 34057 21975 34115 21981
rect 30322 21916 32168 21944
rect 32324 21916 33180 21944
rect 33229 21947 33287 21953
rect 30322 21913 30334 21916
rect 30276 21907 30334 21913
rect 31386 21876 31392 21888
rect 27540 21848 31392 21876
rect 31386 21836 31392 21848
rect 31444 21836 31450 21888
rect 32140 21885 32168 21916
rect 33229 21913 33241 21947
rect 33275 21944 33287 21947
rect 33502 21944 33508 21956
rect 33275 21916 33508 21944
rect 33275 21913 33287 21916
rect 33229 21907 33287 21913
rect 33502 21904 33508 21916
rect 33560 21904 33566 21956
rect 34072 21944 34100 21975
rect 34146 21972 34152 22024
rect 34204 22012 34210 22024
rect 35253 22015 35311 22021
rect 34204 21984 34297 22012
rect 34204 21972 34210 21984
rect 35253 21981 35265 22015
rect 35299 22012 35311 22015
rect 35894 22012 35900 22024
rect 35299 21984 35900 22012
rect 35299 21981 35311 21984
rect 35253 21975 35311 21981
rect 35894 21972 35900 21984
rect 35952 21972 35958 22024
rect 36004 22012 36032 22052
rect 36170 22040 36176 22052
rect 36228 22040 36234 22092
rect 36262 22012 36268 22024
rect 36004 21984 36268 22012
rect 36262 21972 36268 21984
rect 36320 21972 36326 22024
rect 37550 22012 37556 22024
rect 37511 21984 37556 22012
rect 37550 21972 37556 21984
rect 37608 21972 37614 22024
rect 35158 21944 35164 21956
rect 34072 21916 35164 21944
rect 35158 21904 35164 21916
rect 35216 21904 35222 21956
rect 35989 21947 36047 21953
rect 35989 21944 36001 21947
rect 35360 21916 36001 21944
rect 35360 21888 35388 21916
rect 35989 21913 36001 21916
rect 36035 21913 36047 21947
rect 35989 21907 36047 21913
rect 32125 21879 32183 21885
rect 32125 21845 32137 21879
rect 32171 21845 32183 21879
rect 35342 21876 35348 21888
rect 35303 21848 35348 21876
rect 32125 21839 32183 21845
rect 35342 21836 35348 21848
rect 35400 21836 35406 21888
rect 35618 21836 35624 21888
rect 35676 21876 35682 21888
rect 36449 21879 36507 21885
rect 36449 21876 36461 21879
rect 35676 21848 36461 21876
rect 35676 21836 35682 21848
rect 36449 21845 36461 21848
rect 36495 21845 36507 21879
rect 36449 21839 36507 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 18877 21675 18935 21681
rect 18877 21641 18889 21675
rect 18923 21672 18935 21675
rect 19058 21672 19064 21684
rect 18923 21644 19064 21672
rect 18923 21641 18935 21644
rect 18877 21635 18935 21641
rect 19058 21632 19064 21644
rect 19116 21632 19122 21684
rect 21174 21672 21180 21684
rect 21135 21644 21180 21672
rect 21174 21632 21180 21644
rect 21232 21632 21238 21684
rect 23198 21632 23204 21684
rect 23256 21672 23262 21684
rect 23385 21675 23443 21681
rect 23385 21672 23397 21675
rect 23256 21644 23397 21672
rect 23256 21632 23262 21644
rect 23385 21641 23397 21644
rect 23431 21641 23443 21675
rect 27982 21672 27988 21684
rect 27943 21644 27988 21672
rect 23385 21635 23443 21641
rect 27982 21632 27988 21644
rect 28040 21632 28046 21684
rect 28534 21632 28540 21684
rect 28592 21672 28598 21684
rect 29365 21675 29423 21681
rect 29365 21672 29377 21675
rect 28592 21644 29377 21672
rect 28592 21632 28598 21644
rect 29365 21641 29377 21644
rect 29411 21641 29423 21675
rect 31754 21672 31760 21684
rect 29365 21635 29423 21641
rect 29932 21644 31760 21672
rect 19812 21576 22048 21604
rect 17862 21496 17868 21548
rect 17920 21536 17926 21548
rect 18601 21539 18659 21545
rect 18601 21536 18613 21539
rect 17920 21508 18613 21536
rect 17920 21496 17926 21508
rect 18601 21505 18613 21508
rect 18647 21505 18659 21539
rect 18601 21499 18659 21505
rect 18693 21539 18751 21545
rect 18693 21505 18705 21539
rect 18739 21536 18751 21539
rect 18782 21536 18788 21548
rect 18739 21508 18788 21536
rect 18739 21505 18751 21508
rect 18693 21499 18751 21505
rect 18782 21496 18788 21508
rect 18840 21496 18846 21548
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19812 21545 19840 21576
rect 22020 21548 22048 21576
rect 22094 21564 22100 21616
rect 22152 21604 22158 21616
rect 22250 21607 22308 21613
rect 22250 21604 22262 21607
rect 22152 21576 22262 21604
rect 22152 21564 22158 21576
rect 22250 21573 22262 21576
rect 22296 21573 22308 21607
rect 27525 21607 27583 21613
rect 27525 21604 27537 21607
rect 22250 21567 22308 21573
rect 26620 21576 27537 21604
rect 19797 21539 19855 21545
rect 19797 21536 19809 21539
rect 19484 21508 19809 21536
rect 19484 21496 19490 21508
rect 19797 21505 19809 21508
rect 19843 21505 19855 21539
rect 19797 21499 19855 21505
rect 19886 21496 19892 21548
rect 19944 21496 19950 21548
rect 20070 21545 20076 21548
rect 20064 21536 20076 21545
rect 20031 21508 20076 21536
rect 20064 21499 20076 21508
rect 20070 21496 20076 21499
rect 20128 21496 20134 21548
rect 22002 21536 22008 21548
rect 21915 21508 22008 21536
rect 22002 21496 22008 21508
rect 22060 21496 22066 21548
rect 23566 21496 23572 21548
rect 23624 21536 23630 21548
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23624 21508 23857 21536
rect 23624 21496 23630 21508
rect 23845 21505 23857 21508
rect 23891 21505 23903 21539
rect 24026 21536 24032 21548
rect 23987 21508 24032 21536
rect 23845 21499 23903 21505
rect 24026 21496 24032 21508
rect 24084 21496 24090 21548
rect 24210 21496 24216 21548
rect 24268 21536 24274 21548
rect 24765 21539 24823 21545
rect 24765 21536 24777 21539
rect 24268 21508 24777 21536
rect 24268 21496 24274 21508
rect 24765 21505 24777 21508
rect 24811 21536 24823 21539
rect 25038 21536 25044 21548
rect 24811 21508 25044 21536
rect 24811 21505 24823 21508
rect 24765 21499 24823 21505
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21536 25927 21539
rect 26234 21536 26240 21548
rect 25915 21508 26240 21536
rect 25915 21505 25927 21508
rect 25869 21499 25927 21505
rect 26234 21496 26240 21508
rect 26292 21496 26298 21548
rect 26620 21545 26648 21576
rect 27525 21573 27537 21576
rect 27571 21573 27583 21607
rect 27525 21567 27583 21573
rect 28184 21576 29224 21604
rect 26605 21539 26663 21545
rect 26605 21505 26617 21539
rect 26651 21505 26663 21539
rect 27338 21536 27344 21548
rect 27299 21508 27344 21536
rect 26605 21499 26663 21505
rect 27338 21496 27344 21508
rect 27396 21536 27402 21548
rect 28184 21536 28212 21576
rect 27396 21508 28212 21536
rect 28261 21539 28319 21545
rect 27396 21496 27402 21508
rect 28261 21505 28273 21539
rect 28307 21536 28319 21539
rect 28810 21536 28816 21548
rect 28307 21508 28816 21536
rect 28307 21505 28319 21508
rect 28261 21499 28319 21505
rect 28810 21496 28816 21508
rect 28868 21496 28874 21548
rect 29196 21545 29224 21576
rect 29932 21548 29960 21644
rect 31754 21632 31760 21644
rect 31812 21632 31818 21684
rect 32309 21675 32367 21681
rect 32309 21641 32321 21675
rect 32355 21672 32367 21675
rect 32582 21672 32588 21684
rect 32355 21644 32588 21672
rect 32355 21641 32367 21644
rect 32309 21635 32367 21641
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 33597 21675 33655 21681
rect 33597 21641 33609 21675
rect 33643 21672 33655 21675
rect 35710 21672 35716 21684
rect 33643 21644 35716 21672
rect 33643 21641 33655 21644
rect 33597 21635 33655 21641
rect 35710 21632 35716 21644
rect 35768 21672 35774 21684
rect 35768 21644 35894 21672
rect 35768 21632 35774 21644
rect 30101 21607 30159 21613
rect 30101 21573 30113 21607
rect 30147 21604 30159 21607
rect 30282 21604 30288 21616
rect 30147 21576 30288 21604
rect 30147 21573 30159 21576
rect 30101 21567 30159 21573
rect 30282 21564 30288 21576
rect 30340 21604 30346 21616
rect 31021 21607 31079 21613
rect 31021 21604 31033 21607
rect 30340 21576 31033 21604
rect 30340 21564 30346 21576
rect 31021 21573 31033 21576
rect 31067 21573 31079 21607
rect 31021 21567 31079 21573
rect 29181 21539 29239 21545
rect 29181 21505 29193 21539
rect 29227 21536 29239 21539
rect 29914 21536 29920 21548
rect 29227 21508 29920 21536
rect 29227 21505 29239 21508
rect 29181 21499 29239 21505
rect 29914 21496 29920 21508
rect 29972 21496 29978 21548
rect 31036 21536 31064 21567
rect 31386 21564 31392 21616
rect 31444 21604 31450 21616
rect 33502 21604 33508 21616
rect 31444 21576 32812 21604
rect 31444 21564 31450 21576
rect 32582 21536 32588 21548
rect 31036 21508 32444 21536
rect 32543 21508 32588 21536
rect 18877 21471 18935 21477
rect 18877 21437 18889 21471
rect 18923 21468 18935 21471
rect 19904 21468 19932 21496
rect 18923 21440 19932 21468
rect 27157 21471 27215 21477
rect 18923 21437 18935 21440
rect 18877 21431 18935 21437
rect 27157 21437 27169 21471
rect 27203 21468 27215 21471
rect 27522 21468 27528 21480
rect 27203 21440 27528 21468
rect 27203 21437 27215 21440
rect 27157 21431 27215 21437
rect 27522 21428 27528 21440
rect 27580 21428 27586 21480
rect 28166 21468 28172 21480
rect 28127 21440 28172 21468
rect 28166 21428 28172 21440
rect 28224 21428 28230 21480
rect 28353 21471 28411 21477
rect 28353 21437 28365 21471
rect 28399 21437 28411 21471
rect 28353 21431 28411 21437
rect 28074 21360 28080 21412
rect 28132 21400 28138 21412
rect 28368 21400 28396 21431
rect 28442 21428 28448 21480
rect 28500 21468 28506 21480
rect 28500 21440 28545 21468
rect 28500 21428 28506 21440
rect 28626 21428 28632 21480
rect 28684 21468 28690 21480
rect 28997 21471 29055 21477
rect 28997 21468 29009 21471
rect 28684 21440 29009 21468
rect 28684 21428 28690 21440
rect 28997 21437 29009 21440
rect 29043 21437 29055 21471
rect 28997 21431 29055 21437
rect 28902 21400 28908 21412
rect 28132 21372 28908 21400
rect 28132 21360 28138 21372
rect 28902 21360 28908 21372
rect 28960 21400 28966 21412
rect 30377 21403 30435 21409
rect 30377 21400 30389 21403
rect 28960 21372 30389 21400
rect 28960 21360 28966 21372
rect 30377 21369 30389 21372
rect 30423 21369 30435 21403
rect 30377 21363 30435 21369
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 23845 21335 23903 21341
rect 23845 21332 23857 21335
rect 23532 21304 23857 21332
rect 23532 21292 23538 21304
rect 23845 21301 23857 21304
rect 23891 21301 23903 21335
rect 23845 21295 23903 21301
rect 25041 21335 25099 21341
rect 25041 21301 25053 21335
rect 25087 21332 25099 21335
rect 25222 21332 25228 21344
rect 25087 21304 25228 21332
rect 25087 21301 25099 21304
rect 25041 21295 25099 21301
rect 25222 21292 25228 21304
rect 25280 21292 25286 21344
rect 25498 21292 25504 21344
rect 25556 21332 25562 21344
rect 25685 21335 25743 21341
rect 25685 21332 25697 21335
rect 25556 21304 25697 21332
rect 25556 21292 25562 21304
rect 25685 21301 25697 21304
rect 25731 21301 25743 21335
rect 25685 21295 25743 21301
rect 26421 21335 26479 21341
rect 26421 21301 26433 21335
rect 26467 21332 26479 21335
rect 26694 21332 26700 21344
rect 26467 21304 26700 21332
rect 26467 21301 26479 21304
rect 26421 21295 26479 21301
rect 26694 21292 26700 21304
rect 26752 21292 26758 21344
rect 30926 21292 30932 21344
rect 30984 21332 30990 21344
rect 31113 21335 31171 21341
rect 31113 21332 31125 21335
rect 30984 21304 31125 21332
rect 30984 21292 30990 21304
rect 31113 21301 31125 21304
rect 31159 21301 31171 21335
rect 32416 21332 32444 21508
rect 32582 21496 32588 21508
rect 32640 21496 32646 21548
rect 32784 21545 32812 21576
rect 32968 21576 33508 21604
rect 32968 21545 32996 21576
rect 33502 21564 33508 21576
rect 33560 21564 33566 21616
rect 34698 21604 34704 21616
rect 34532 21576 34704 21604
rect 34532 21545 34560 21576
rect 34698 21564 34704 21576
rect 34756 21564 34762 21616
rect 34793 21607 34851 21613
rect 34793 21573 34805 21607
rect 34839 21604 34851 21607
rect 35618 21604 35624 21616
rect 34839 21576 35624 21604
rect 34839 21573 34851 21576
rect 34793 21567 34851 21573
rect 35618 21564 35624 21576
rect 35676 21564 35682 21616
rect 35866 21604 35894 21644
rect 36170 21632 36176 21684
rect 36228 21672 36234 21684
rect 36633 21675 36691 21681
rect 36633 21672 36645 21675
rect 36228 21644 36645 21672
rect 36228 21632 36234 21644
rect 36633 21641 36645 21644
rect 36679 21641 36691 21675
rect 36633 21635 36691 21641
rect 37642 21604 37648 21616
rect 35866 21576 37648 21604
rect 37642 21564 37648 21576
rect 37700 21564 37706 21616
rect 32677 21539 32735 21545
rect 32677 21505 32689 21539
rect 32723 21505 32735 21539
rect 32677 21499 32735 21505
rect 32769 21539 32827 21545
rect 32769 21505 32781 21539
rect 32815 21505 32827 21539
rect 32769 21499 32827 21505
rect 32953 21539 33011 21545
rect 32953 21505 32965 21539
rect 32999 21505 33011 21539
rect 32953 21499 33011 21505
rect 34517 21539 34575 21545
rect 34517 21505 34529 21539
rect 34563 21505 34575 21539
rect 34517 21499 34575 21505
rect 34609 21539 34667 21545
rect 34609 21505 34621 21539
rect 34655 21505 34667 21539
rect 34609 21499 34667 21505
rect 35520 21539 35578 21545
rect 35520 21505 35532 21539
rect 35566 21536 35578 21539
rect 36630 21536 36636 21548
rect 35566 21508 36636 21536
rect 35566 21505 35578 21508
rect 35520 21499 35578 21505
rect 32692 21412 32720 21499
rect 32674 21360 32680 21412
rect 32732 21360 32738 21412
rect 32968 21332 32996 21499
rect 34146 21428 34152 21480
rect 34204 21468 34210 21480
rect 34624 21468 34652 21499
rect 36630 21496 36636 21508
rect 36688 21496 36694 21548
rect 34790 21468 34796 21480
rect 34204 21440 34796 21468
rect 34204 21428 34210 21440
rect 34790 21428 34796 21440
rect 34848 21428 34854 21480
rect 35253 21471 35311 21477
rect 35253 21437 35265 21471
rect 35299 21437 35311 21471
rect 35253 21431 35311 21437
rect 32416 21304 32996 21332
rect 35268 21332 35296 21431
rect 35526 21332 35532 21344
rect 35268 21304 35532 21332
rect 31113 21295 31171 21301
rect 35526 21292 35532 21304
rect 35584 21292 35590 21344
rect 35618 21292 35624 21344
rect 35676 21332 35682 21344
rect 36170 21332 36176 21344
rect 35676 21304 36176 21332
rect 35676 21292 35682 21304
rect 36170 21292 36176 21304
rect 36228 21292 36234 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 23566 21088 23572 21140
rect 23624 21128 23630 21140
rect 23845 21131 23903 21137
rect 23845 21128 23857 21131
rect 23624 21100 23857 21128
rect 23624 21088 23630 21100
rect 23845 21097 23857 21100
rect 23891 21097 23903 21131
rect 23845 21091 23903 21097
rect 28166 21088 28172 21140
rect 28224 21128 28230 21140
rect 28813 21131 28871 21137
rect 28813 21128 28825 21131
rect 28224 21100 28825 21128
rect 28224 21088 28230 21100
rect 28813 21097 28825 21100
rect 28859 21097 28871 21131
rect 28813 21091 28871 21097
rect 27801 21063 27859 21069
rect 27801 21029 27813 21063
rect 27847 21060 27859 21063
rect 28350 21060 28356 21072
rect 27847 21032 28356 21060
rect 27847 21029 27859 21032
rect 27801 21023 27859 21029
rect 28350 21020 28356 21032
rect 28408 21060 28414 21072
rect 28626 21060 28632 21072
rect 28408 21032 28632 21060
rect 28408 21020 28414 21032
rect 28626 21020 28632 21032
rect 28684 21020 28690 21072
rect 24302 20952 24308 21004
rect 24360 20992 24366 21004
rect 24581 20995 24639 21001
rect 24581 20992 24593 20995
rect 24360 20964 24593 20992
rect 24360 20952 24366 20964
rect 24581 20961 24593 20964
rect 24627 20961 24639 20995
rect 24581 20955 24639 20961
rect 29730 20952 29736 21004
rect 29788 20992 29794 21004
rect 30006 20992 30012 21004
rect 29788 20964 30012 20992
rect 29788 20952 29794 20964
rect 30006 20952 30012 20964
rect 30064 20992 30070 21004
rect 30285 20995 30343 21001
rect 30285 20992 30297 20995
rect 30064 20964 30297 20992
rect 30064 20952 30070 20964
rect 30285 20961 30297 20964
rect 30331 20961 30343 20995
rect 30285 20955 30343 20961
rect 1762 20924 1768 20936
rect 1723 20896 1768 20924
rect 1762 20884 1768 20896
rect 1820 20884 1826 20936
rect 22002 20884 22008 20936
rect 22060 20924 22066 20936
rect 22465 20927 22523 20933
rect 22465 20924 22477 20927
rect 22060 20896 22477 20924
rect 22060 20884 22066 20896
rect 22465 20893 22477 20896
rect 22511 20924 22523 20927
rect 23566 20924 23572 20936
rect 22511 20896 23572 20924
rect 22511 20893 22523 20896
rect 22465 20887 22523 20893
rect 23566 20884 23572 20896
rect 23624 20924 23630 20936
rect 24320 20924 24348 20952
rect 23624 20896 24348 20924
rect 26421 20927 26479 20933
rect 23624 20884 23630 20896
rect 26421 20893 26433 20927
rect 26467 20924 26479 20927
rect 27706 20924 27712 20936
rect 26467 20896 27712 20924
rect 26467 20893 26479 20896
rect 26421 20887 26479 20893
rect 27706 20884 27712 20896
rect 27764 20884 27770 20936
rect 28626 20924 28632 20936
rect 28587 20896 28632 20924
rect 28626 20884 28632 20896
rect 28684 20884 28690 20936
rect 30558 20933 30564 20936
rect 30552 20887 30564 20933
rect 30616 20924 30622 20936
rect 30616 20896 30652 20924
rect 30558 20884 30564 20887
rect 30616 20884 30622 20896
rect 32398 20884 32404 20936
rect 32456 20924 32462 20936
rect 32677 20927 32735 20933
rect 32677 20924 32689 20927
rect 32456 20896 32689 20924
rect 32456 20884 32462 20896
rect 32677 20893 32689 20896
rect 32723 20893 32735 20927
rect 32677 20887 32735 20893
rect 34885 20927 34943 20933
rect 34885 20893 34897 20927
rect 34931 20924 34943 20927
rect 35526 20924 35532 20936
rect 34931 20896 35532 20924
rect 34931 20893 34943 20896
rect 34885 20887 34943 20893
rect 35526 20884 35532 20896
rect 35584 20884 35590 20936
rect 22732 20859 22790 20865
rect 22732 20825 22744 20859
rect 22778 20856 22790 20859
rect 23474 20856 23480 20868
rect 22778 20828 23480 20856
rect 22778 20825 22790 20828
rect 22732 20819 22790 20825
rect 23474 20816 23480 20828
rect 23532 20816 23538 20868
rect 24854 20865 24860 20868
rect 24848 20819 24860 20865
rect 24912 20856 24918 20868
rect 26694 20865 26700 20868
rect 26688 20856 26700 20865
rect 24912 20828 24948 20856
rect 26655 20828 26700 20856
rect 24854 20816 24860 20819
rect 24912 20816 24918 20828
rect 26688 20819 26700 20828
rect 26694 20816 26700 20819
rect 26752 20816 26758 20868
rect 27522 20816 27528 20868
rect 27580 20856 27586 20868
rect 28261 20859 28319 20865
rect 28261 20856 28273 20859
rect 27580 20828 28273 20856
rect 27580 20816 27586 20828
rect 28261 20825 28273 20828
rect 28307 20825 28319 20859
rect 28261 20819 28319 20825
rect 32944 20859 33002 20865
rect 32944 20825 32956 20859
rect 32990 20856 33002 20859
rect 33134 20856 33140 20868
rect 32990 20828 33140 20856
rect 32990 20825 33002 20828
rect 32944 20819 33002 20825
rect 33134 20816 33140 20828
rect 33192 20816 33198 20868
rect 35152 20859 35210 20865
rect 35152 20825 35164 20859
rect 35198 20856 35210 20859
rect 35986 20856 35992 20868
rect 35198 20828 35992 20856
rect 35198 20825 35210 20828
rect 35152 20819 35210 20825
rect 35986 20816 35992 20828
rect 36044 20816 36050 20868
rect 25130 20748 25136 20800
rect 25188 20788 25194 20800
rect 25961 20791 26019 20797
rect 25961 20788 25973 20791
rect 25188 20760 25973 20788
rect 25188 20748 25194 20760
rect 25961 20757 25973 20760
rect 26007 20757 26019 20791
rect 25961 20751 26019 20757
rect 27982 20748 27988 20800
rect 28040 20788 28046 20800
rect 28445 20791 28503 20797
rect 28445 20788 28457 20791
rect 28040 20760 28457 20788
rect 28040 20748 28046 20760
rect 28445 20757 28457 20760
rect 28491 20757 28503 20791
rect 28445 20751 28503 20757
rect 28534 20748 28540 20800
rect 28592 20788 28598 20800
rect 31662 20788 31668 20800
rect 28592 20760 28637 20788
rect 31623 20760 31668 20788
rect 28592 20748 28598 20760
rect 31662 20748 31668 20760
rect 31720 20748 31726 20800
rect 32490 20748 32496 20800
rect 32548 20788 32554 20800
rect 34057 20791 34115 20797
rect 34057 20788 34069 20791
rect 32548 20760 34069 20788
rect 32548 20748 32554 20760
rect 34057 20757 34069 20760
rect 34103 20757 34115 20791
rect 34057 20751 34115 20757
rect 35250 20748 35256 20800
rect 35308 20788 35314 20800
rect 36265 20791 36323 20797
rect 36265 20788 36277 20791
rect 35308 20760 36277 20788
rect 35308 20748 35314 20760
rect 36265 20757 36277 20760
rect 36311 20757 36323 20791
rect 36265 20751 36323 20757
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 24397 20587 24455 20593
rect 24397 20553 24409 20587
rect 24443 20584 24455 20587
rect 24854 20584 24860 20596
rect 24443 20556 24860 20584
rect 24443 20553 24455 20556
rect 24397 20547 24455 20553
rect 24854 20544 24860 20556
rect 24912 20544 24918 20596
rect 29086 20584 29092 20596
rect 28184 20556 29092 20584
rect 19705 20519 19763 20525
rect 19705 20485 19717 20519
rect 19751 20516 19763 20519
rect 19751 20488 20760 20516
rect 19751 20485 19763 20488
rect 19705 20479 19763 20485
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20448 20591 20451
rect 20622 20448 20628 20460
rect 20579 20420 20628 20448
rect 20579 20417 20591 20420
rect 20533 20411 20591 20417
rect 20622 20408 20628 20420
rect 20680 20408 20686 20460
rect 20732 20457 20760 20488
rect 24026 20476 24032 20528
rect 24084 20516 24090 20528
rect 27706 20516 27712 20528
rect 24084 20488 24532 20516
rect 24084 20476 24090 20488
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20448 20775 20451
rect 24210 20448 24216 20460
rect 20763 20420 24216 20448
rect 20763 20417 20775 20420
rect 20717 20411 20775 20417
rect 24210 20408 24216 20420
rect 24268 20408 24274 20460
rect 24504 20457 24532 20488
rect 25240 20488 27712 20516
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 24489 20451 24547 20457
rect 24489 20417 24501 20451
rect 24535 20448 24547 20451
rect 24854 20448 24860 20460
rect 24535 20420 24860 20448
rect 24535 20417 24547 20420
rect 24489 20411 24547 20417
rect 24320 20380 24348 20411
rect 24854 20408 24860 20420
rect 24912 20408 24918 20460
rect 25240 20457 25268 20488
rect 27706 20476 27712 20488
rect 27764 20476 27770 20528
rect 25498 20457 25504 20460
rect 25225 20451 25283 20457
rect 25225 20417 25237 20451
rect 25271 20417 25283 20451
rect 25492 20448 25504 20457
rect 25459 20420 25504 20448
rect 25225 20411 25283 20417
rect 25492 20411 25504 20420
rect 25498 20408 25504 20411
rect 25556 20408 25562 20460
rect 27522 20448 27528 20460
rect 26620 20420 27528 20448
rect 25130 20380 25136 20392
rect 24320 20352 25136 20380
rect 25130 20340 25136 20352
rect 25188 20340 25194 20392
rect 24026 20312 24032 20324
rect 20088 20284 24032 20312
rect 20088 20256 20116 20284
rect 24026 20272 24032 20284
rect 24084 20272 24090 20324
rect 26620 20321 26648 20420
rect 27522 20408 27528 20420
rect 27580 20448 27586 20460
rect 27893 20451 27951 20457
rect 27893 20448 27905 20451
rect 27580 20420 27905 20448
rect 27580 20408 27586 20420
rect 27893 20417 27905 20420
rect 27939 20417 27951 20451
rect 27893 20411 27951 20417
rect 27982 20408 27988 20460
rect 28040 20448 28046 20460
rect 28184 20457 28212 20556
rect 29086 20544 29092 20556
rect 29144 20544 29150 20596
rect 31110 20544 31116 20596
rect 31168 20584 31174 20596
rect 31297 20587 31355 20593
rect 31297 20584 31309 20587
rect 31168 20556 31309 20584
rect 31168 20544 31174 20556
rect 31297 20553 31309 20556
rect 31343 20553 31355 20587
rect 31297 20547 31355 20553
rect 32582 20544 32588 20596
rect 32640 20584 32646 20596
rect 32769 20587 32827 20593
rect 32769 20584 32781 20587
rect 32640 20556 32781 20584
rect 32640 20544 32646 20556
rect 32769 20553 32781 20556
rect 32815 20553 32827 20587
rect 32769 20547 32827 20553
rect 33134 20544 33140 20596
rect 33192 20584 33198 20596
rect 34057 20587 34115 20593
rect 34057 20584 34069 20587
rect 33192 20556 34069 20584
rect 33192 20544 33198 20556
rect 34057 20553 34069 20556
rect 34103 20553 34115 20587
rect 35986 20584 35992 20596
rect 35947 20556 35992 20584
rect 34057 20547 34115 20553
rect 35986 20544 35992 20556
rect 36044 20544 36050 20596
rect 36630 20584 36636 20596
rect 36591 20556 36636 20584
rect 36630 20544 36636 20556
rect 36688 20544 36694 20596
rect 28994 20525 29000 20528
rect 28988 20479 29000 20525
rect 29052 20516 29058 20528
rect 32309 20519 32367 20525
rect 32309 20516 32321 20519
rect 29052 20488 29088 20516
rect 31036 20488 32321 20516
rect 28994 20476 29000 20479
rect 29052 20476 29058 20488
rect 31036 20457 31064 20488
rect 32309 20485 32321 20488
rect 32355 20516 32367 20519
rect 32490 20516 32496 20528
rect 32355 20488 32496 20516
rect 32355 20485 32367 20488
rect 32309 20479 32367 20485
rect 32490 20476 32496 20488
rect 32548 20476 32554 20528
rect 34790 20476 34796 20528
rect 34848 20516 34854 20528
rect 35529 20519 35587 20525
rect 34848 20488 35388 20516
rect 34848 20476 34854 20488
rect 28169 20451 28227 20457
rect 28040 20420 28085 20448
rect 28040 20408 28046 20420
rect 28169 20417 28181 20451
rect 28215 20417 28227 20451
rect 28169 20411 28227 20417
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20417 31079 20451
rect 31021 20411 31079 20417
rect 31113 20451 31171 20457
rect 31113 20417 31125 20451
rect 31159 20417 31171 20451
rect 31113 20411 31171 20417
rect 32585 20451 32643 20457
rect 32585 20417 32597 20451
rect 32631 20417 32643 20451
rect 32585 20411 32643 20417
rect 33413 20451 33471 20457
rect 33413 20417 33425 20451
rect 33459 20448 33471 20451
rect 33502 20448 33508 20460
rect 33459 20420 33508 20448
rect 33459 20417 33471 20420
rect 33413 20411 33471 20417
rect 27706 20340 27712 20392
rect 27764 20380 27770 20392
rect 28721 20383 28779 20389
rect 28721 20380 28733 20383
rect 27764 20352 28733 20380
rect 27764 20340 27770 20352
rect 28721 20349 28733 20352
rect 28767 20349 28779 20383
rect 28721 20343 28779 20349
rect 30558 20340 30564 20392
rect 30616 20380 30622 20392
rect 30926 20380 30932 20392
rect 30616 20352 30932 20380
rect 30616 20340 30622 20352
rect 30926 20340 30932 20352
rect 30984 20380 30990 20392
rect 31128 20380 31156 20411
rect 30984 20352 31156 20380
rect 30984 20340 30990 20352
rect 31662 20340 31668 20392
rect 31720 20380 31726 20392
rect 32493 20383 32551 20389
rect 32493 20380 32505 20383
rect 31720 20352 32505 20380
rect 31720 20340 31726 20352
rect 32493 20349 32505 20352
rect 32539 20349 32551 20383
rect 32600 20380 32628 20411
rect 33502 20408 33508 20420
rect 33560 20408 33566 20460
rect 33597 20451 33655 20457
rect 33597 20417 33609 20451
rect 33643 20448 33655 20451
rect 34241 20451 34299 20457
rect 34241 20448 34253 20451
rect 33643 20420 34253 20448
rect 33643 20417 33655 20420
rect 33597 20411 33655 20417
rect 34241 20417 34253 20420
rect 34287 20417 34299 20451
rect 35250 20448 35256 20460
rect 35211 20420 35256 20448
rect 34241 20411 34299 20417
rect 35250 20408 35256 20420
rect 35308 20408 35314 20460
rect 35360 20457 35388 20488
rect 35529 20485 35541 20519
rect 35575 20516 35587 20519
rect 35575 20488 36860 20516
rect 35575 20485 35587 20488
rect 35529 20479 35587 20485
rect 35345 20451 35403 20457
rect 35345 20417 35357 20451
rect 35391 20417 35403 20451
rect 36170 20448 36176 20460
rect 36131 20420 36176 20448
rect 35345 20411 35403 20417
rect 36170 20408 36176 20420
rect 36228 20408 36234 20460
rect 36832 20457 36860 20488
rect 36817 20451 36875 20457
rect 36817 20417 36829 20451
rect 36863 20417 36875 20451
rect 36817 20411 36875 20417
rect 33226 20380 33232 20392
rect 32600 20352 33232 20380
rect 32493 20343 32551 20349
rect 26605 20315 26663 20321
rect 26605 20281 26617 20315
rect 26651 20281 26663 20315
rect 26605 20275 26663 20281
rect 28077 20315 28135 20321
rect 28077 20281 28089 20315
rect 28123 20312 28135 20315
rect 28626 20312 28632 20324
rect 28123 20284 28632 20312
rect 28123 20281 28135 20284
rect 28077 20275 28135 20281
rect 28626 20272 28632 20284
rect 28684 20272 28690 20324
rect 32508 20312 32536 20343
rect 33226 20340 33232 20352
rect 33284 20340 33290 20392
rect 33318 20312 33324 20324
rect 32508 20284 33324 20312
rect 33318 20272 33324 20284
rect 33376 20272 33382 20324
rect 19981 20247 20039 20253
rect 19981 20213 19993 20247
rect 20027 20244 20039 20247
rect 20070 20244 20076 20256
rect 20027 20216 20076 20244
rect 20027 20213 20039 20216
rect 19981 20207 20039 20213
rect 20070 20204 20076 20216
rect 20128 20204 20134 20256
rect 20530 20244 20536 20256
rect 20491 20216 20536 20244
rect 20530 20204 20536 20216
rect 20588 20204 20594 20256
rect 27709 20247 27767 20253
rect 27709 20213 27721 20247
rect 27755 20244 27767 20247
rect 28442 20244 28448 20256
rect 27755 20216 28448 20244
rect 27755 20213 27767 20216
rect 27709 20207 27767 20213
rect 28442 20204 28448 20216
rect 28500 20204 28506 20256
rect 28534 20204 28540 20256
rect 28592 20244 28598 20256
rect 30101 20247 30159 20253
rect 30101 20244 30113 20247
rect 28592 20216 30113 20244
rect 28592 20204 28598 20216
rect 30101 20213 30113 20216
rect 30147 20213 30159 20247
rect 30101 20207 30159 20213
rect 31386 20204 31392 20256
rect 31444 20244 31450 20256
rect 32309 20247 32367 20253
rect 32309 20244 32321 20247
rect 31444 20216 32321 20244
rect 31444 20204 31450 20216
rect 32309 20213 32321 20216
rect 32355 20244 32367 20247
rect 33134 20244 33140 20256
rect 32355 20216 33140 20244
rect 32355 20213 32367 20216
rect 32309 20207 32367 20213
rect 33134 20204 33140 20216
rect 33192 20204 33198 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 26234 20040 26240 20052
rect 26195 20012 26240 20040
rect 26234 20000 26240 20012
rect 26292 20000 26298 20052
rect 28350 20040 28356 20052
rect 28311 20012 28356 20040
rect 28350 20000 28356 20012
rect 28408 20000 28414 20052
rect 28626 20040 28632 20052
rect 28587 20012 28632 20040
rect 28626 20000 28632 20012
rect 28684 20000 28690 20052
rect 33226 20000 33232 20052
rect 33284 20040 33290 20052
rect 33873 20043 33931 20049
rect 33873 20040 33885 20043
rect 33284 20012 33885 20040
rect 33284 20000 33290 20012
rect 33873 20009 33885 20012
rect 33919 20009 33931 20043
rect 33873 20003 33931 20009
rect 24857 19975 24915 19981
rect 24857 19941 24869 19975
rect 24903 19972 24915 19975
rect 25774 19972 25780 19984
rect 24903 19944 25780 19972
rect 24903 19941 24915 19944
rect 24857 19935 24915 19941
rect 25774 19932 25780 19944
rect 25832 19932 25838 19984
rect 25590 19864 25596 19916
rect 25648 19904 25654 19916
rect 25869 19907 25927 19913
rect 25869 19904 25881 19907
rect 25648 19876 25881 19904
rect 25648 19864 25654 19876
rect 25869 19873 25881 19876
rect 25915 19904 25927 19907
rect 27982 19904 27988 19916
rect 25915 19876 27988 19904
rect 25915 19873 25927 19876
rect 25869 19867 25927 19873
rect 27982 19864 27988 19876
rect 28040 19864 28046 19916
rect 31113 19907 31171 19913
rect 31113 19873 31125 19907
rect 31159 19904 31171 19907
rect 31662 19904 31668 19916
rect 31159 19876 31668 19904
rect 31159 19873 31171 19876
rect 31113 19867 31171 19873
rect 31662 19864 31668 19876
rect 31720 19864 31726 19916
rect 33502 19864 33508 19916
rect 33560 19904 33566 19916
rect 33560 19876 35112 19904
rect 33560 19864 33566 19876
rect 19426 19796 19432 19848
rect 19484 19836 19490 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 19484 19808 19901 19836
rect 19484 19796 19490 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 22186 19836 22192 19848
rect 22147 19808 22192 19836
rect 19889 19799 19947 19805
rect 22186 19796 22192 19808
rect 22244 19796 22250 19848
rect 22373 19839 22431 19845
rect 22373 19805 22385 19839
rect 22419 19805 22431 19839
rect 23842 19836 23848 19848
rect 23803 19808 23848 19836
rect 22373 19799 22431 19805
rect 20156 19771 20214 19777
rect 20156 19737 20168 19771
rect 20202 19768 20214 19771
rect 20346 19768 20352 19780
rect 20202 19740 20352 19768
rect 20202 19737 20214 19740
rect 20156 19731 20214 19737
rect 20346 19728 20352 19740
rect 20404 19728 20410 19780
rect 21634 19728 21640 19780
rect 21692 19768 21698 19780
rect 22388 19768 22416 19799
rect 23842 19796 23848 19808
rect 23900 19796 23906 19848
rect 24026 19836 24032 19848
rect 23987 19808 24032 19836
rect 24026 19796 24032 19808
rect 24084 19796 24090 19848
rect 25130 19836 25136 19848
rect 25091 19808 25136 19836
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 26053 19839 26111 19845
rect 26053 19805 26065 19839
rect 26099 19836 26111 19839
rect 27338 19836 27344 19848
rect 26099 19808 27344 19836
rect 26099 19805 26111 19808
rect 26053 19799 26111 19805
rect 27338 19796 27344 19808
rect 27396 19796 27402 19848
rect 28258 19836 28264 19848
rect 28219 19808 28264 19836
rect 28258 19796 28264 19808
rect 28316 19796 28322 19848
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19836 28503 19839
rect 28534 19836 28540 19848
rect 28491 19808 28540 19836
rect 28491 19805 28503 19808
rect 28445 19799 28503 19805
rect 28534 19796 28540 19808
rect 28592 19836 28598 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 28592 19808 29745 19836
rect 28592 19796 28598 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29914 19836 29920 19848
rect 29875 19808 29920 19836
rect 29733 19799 29791 19805
rect 29914 19796 29920 19808
rect 29972 19796 29978 19848
rect 30558 19796 30564 19848
rect 30616 19836 30622 19848
rect 31297 19839 31355 19845
rect 31297 19836 31309 19839
rect 30616 19808 31309 19836
rect 30616 19796 30622 19808
rect 31297 19805 31309 19808
rect 31343 19836 31355 19839
rect 31570 19836 31576 19848
rect 31343 19808 31576 19836
rect 31343 19805 31355 19808
rect 31297 19799 31355 19805
rect 31570 19796 31576 19808
rect 31628 19796 31634 19848
rect 32398 19796 32404 19848
rect 32456 19836 32462 19848
rect 35084 19845 35112 19876
rect 32493 19839 32551 19845
rect 32493 19836 32505 19839
rect 32456 19808 32505 19836
rect 32456 19796 32462 19808
rect 32493 19805 32505 19808
rect 32539 19805 32551 19839
rect 32493 19799 32551 19805
rect 34977 19839 35035 19845
rect 34977 19805 34989 19839
rect 35023 19805 35035 19839
rect 34977 19799 35035 19805
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19805 35127 19839
rect 35986 19836 35992 19848
rect 35947 19808 35992 19836
rect 35069 19799 35127 19805
rect 21692 19740 22416 19768
rect 24857 19771 24915 19777
rect 21692 19728 21698 19740
rect 24857 19737 24869 19771
rect 24903 19768 24915 19771
rect 25222 19768 25228 19780
rect 24903 19740 25228 19768
rect 24903 19737 24915 19740
rect 24857 19731 24915 19737
rect 25222 19728 25228 19740
rect 25280 19768 25286 19780
rect 27154 19768 27160 19780
rect 25280 19740 27160 19768
rect 25280 19728 25286 19740
rect 27154 19728 27160 19740
rect 27212 19728 27218 19780
rect 32760 19771 32818 19777
rect 32760 19737 32772 19771
rect 32806 19768 32818 19771
rect 33410 19768 33416 19780
rect 32806 19740 33416 19768
rect 32806 19737 32818 19740
rect 32760 19731 32818 19737
rect 33410 19728 33416 19740
rect 33468 19728 33474 19780
rect 34992 19768 35020 19799
rect 35986 19796 35992 19808
rect 36044 19796 36050 19848
rect 36538 19768 36544 19780
rect 34992 19740 36544 19768
rect 36538 19728 36544 19740
rect 36596 19728 36602 19780
rect 21266 19700 21272 19712
rect 21227 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 22278 19700 22284 19712
rect 22239 19672 22284 19700
rect 22278 19660 22284 19672
rect 22336 19660 22342 19712
rect 23474 19660 23480 19712
rect 23532 19700 23538 19712
rect 23937 19703 23995 19709
rect 23937 19700 23949 19703
rect 23532 19672 23949 19700
rect 23532 19660 23538 19672
rect 23937 19669 23949 19672
rect 23983 19669 23995 19703
rect 23937 19663 23995 19669
rect 25041 19703 25099 19709
rect 25041 19669 25053 19703
rect 25087 19700 25099 19703
rect 25958 19700 25964 19712
rect 25087 19672 25964 19700
rect 25087 19669 25099 19672
rect 25041 19663 25099 19669
rect 25958 19660 25964 19672
rect 26016 19660 26022 19712
rect 29454 19660 29460 19712
rect 29512 19700 29518 19712
rect 30101 19703 30159 19709
rect 30101 19700 30113 19703
rect 29512 19672 30113 19700
rect 29512 19660 29518 19672
rect 30101 19669 30113 19672
rect 30147 19669 30159 19703
rect 30101 19663 30159 19669
rect 30926 19660 30932 19712
rect 30984 19700 30990 19712
rect 31481 19703 31539 19709
rect 31481 19700 31493 19703
rect 30984 19672 31493 19700
rect 30984 19660 30990 19672
rect 31481 19669 31493 19672
rect 31527 19669 31539 19703
rect 31481 19663 31539 19669
rect 34698 19660 34704 19712
rect 34756 19700 34762 19712
rect 35253 19703 35311 19709
rect 35253 19700 35265 19703
rect 34756 19672 35265 19700
rect 34756 19660 34762 19672
rect 35253 19669 35265 19672
rect 35299 19669 35311 19703
rect 35802 19700 35808 19712
rect 35763 19672 35808 19700
rect 35253 19663 35311 19669
rect 35802 19660 35808 19672
rect 35860 19660 35866 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 20346 19496 20352 19508
rect 20307 19468 20352 19496
rect 20346 19456 20352 19468
rect 20404 19456 20410 19508
rect 25590 19496 25596 19508
rect 25551 19468 25596 19496
rect 25590 19456 25596 19468
rect 25648 19456 25654 19508
rect 26053 19499 26111 19505
rect 26053 19465 26065 19499
rect 26099 19465 26111 19499
rect 26053 19459 26111 19465
rect 19426 19388 19432 19440
rect 19484 19428 19490 19440
rect 22278 19437 22284 19440
rect 22272 19428 22284 19437
rect 19484 19400 22048 19428
rect 22239 19400 22284 19428
rect 19484 19388 19490 19400
rect 22020 19372 22048 19400
rect 22272 19391 22284 19400
rect 22278 19388 22284 19391
rect 22336 19388 22342 19440
rect 24480 19431 24538 19437
rect 24480 19397 24492 19431
rect 24526 19428 24538 19431
rect 26068 19428 26096 19459
rect 28258 19456 28264 19508
rect 28316 19496 28322 19508
rect 28629 19499 28687 19505
rect 28629 19496 28641 19499
rect 28316 19468 28641 19496
rect 28316 19456 28322 19468
rect 28629 19465 28641 19468
rect 28675 19465 28687 19499
rect 28629 19459 28687 19465
rect 30466 19456 30472 19508
rect 30524 19496 30530 19508
rect 30745 19499 30803 19505
rect 30745 19496 30757 19499
rect 30524 19468 30757 19496
rect 30524 19456 30530 19468
rect 30745 19465 30757 19468
rect 30791 19465 30803 19499
rect 30745 19459 30803 19465
rect 32674 19456 32680 19508
rect 32732 19496 32738 19508
rect 32769 19499 32827 19505
rect 32769 19496 32781 19499
rect 32732 19468 32781 19496
rect 32732 19456 32738 19468
rect 32769 19465 32781 19468
rect 32815 19465 32827 19499
rect 32769 19459 32827 19465
rect 32858 19456 32864 19508
rect 32916 19496 32922 19508
rect 33429 19499 33487 19505
rect 33429 19496 33441 19499
rect 32916 19468 33441 19496
rect 32916 19456 32922 19468
rect 33429 19465 33441 19468
rect 33475 19465 33487 19499
rect 33594 19496 33600 19508
rect 33555 19468 33600 19496
rect 33429 19459 33487 19465
rect 33594 19456 33600 19468
rect 33652 19456 33658 19508
rect 36998 19456 37004 19508
rect 37056 19496 37062 19508
rect 37461 19499 37519 19505
rect 37461 19496 37473 19499
rect 37056 19468 37473 19496
rect 37056 19456 37062 19468
rect 37461 19465 37473 19468
rect 37507 19465 37519 19499
rect 37461 19459 37519 19465
rect 24526 19400 26096 19428
rect 31757 19431 31815 19437
rect 24526 19397 24538 19400
rect 24480 19391 24538 19397
rect 31757 19397 31769 19431
rect 31803 19428 31815 19431
rect 33134 19428 33140 19440
rect 31803 19400 33140 19428
rect 31803 19397 31815 19400
rect 31757 19391 31815 19397
rect 33134 19388 33140 19400
rect 33192 19388 33198 19440
rect 33226 19388 33232 19440
rect 33284 19428 33290 19440
rect 35802 19437 35808 19440
rect 35796 19428 35808 19437
rect 33284 19400 33329 19428
rect 35763 19400 35808 19428
rect 33284 19388 33290 19400
rect 35796 19391 35808 19400
rect 35802 19388 35808 19391
rect 35860 19388 35866 19440
rect 19705 19363 19763 19369
rect 19705 19329 19717 19363
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19360 19947 19363
rect 20530 19360 20536 19372
rect 19935 19332 20392 19360
rect 20491 19332 20536 19360
rect 19935 19329 19947 19332
rect 19889 19323 19947 19329
rect 19720 19292 19748 19323
rect 20162 19292 20168 19304
rect 19720 19264 20168 19292
rect 20162 19252 20168 19264
rect 20220 19252 20226 19304
rect 20364 19292 20392 19332
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 22002 19360 22008 19372
rect 21915 19332 22008 19360
rect 22002 19320 22008 19332
rect 22060 19320 22066 19372
rect 26234 19360 26240 19372
rect 26195 19332 26240 19360
rect 26234 19320 26240 19332
rect 26292 19320 26298 19372
rect 27338 19360 27344 19372
rect 27299 19332 27344 19360
rect 27338 19320 27344 19332
rect 27396 19320 27402 19372
rect 28166 19360 28172 19372
rect 28127 19332 28172 19360
rect 28166 19320 28172 19332
rect 28224 19320 28230 19372
rect 28258 19320 28264 19372
rect 28316 19360 28322 19372
rect 28445 19363 28503 19369
rect 28445 19360 28457 19363
rect 28316 19332 28457 19360
rect 28316 19320 28322 19332
rect 28445 19329 28457 19332
rect 28491 19329 28503 19363
rect 29454 19360 29460 19372
rect 29415 19332 29460 19360
rect 28445 19323 28503 19329
rect 29454 19320 29460 19332
rect 29512 19320 29518 19372
rect 29638 19320 29644 19372
rect 29696 19360 29702 19372
rect 30101 19363 30159 19369
rect 30101 19360 30113 19363
rect 29696 19332 30113 19360
rect 29696 19320 29702 19332
rect 30101 19329 30113 19332
rect 30147 19329 30159 19363
rect 30926 19360 30932 19372
rect 30887 19332 30932 19360
rect 30101 19323 30159 19329
rect 30926 19320 30932 19332
rect 30984 19320 30990 19372
rect 31570 19360 31576 19372
rect 31531 19332 31576 19360
rect 31570 19320 31576 19332
rect 31628 19320 31634 19372
rect 32306 19360 32312 19372
rect 32267 19332 32312 19360
rect 32306 19320 32312 19332
rect 32364 19320 32370 19372
rect 32582 19360 32588 19372
rect 32543 19332 32588 19360
rect 32582 19320 32588 19332
rect 32640 19320 32646 19372
rect 34698 19360 34704 19372
rect 34659 19332 34704 19360
rect 34698 19320 34704 19332
rect 34756 19320 34762 19372
rect 37642 19360 37648 19372
rect 37603 19332 37648 19360
rect 37642 19320 37648 19332
rect 37700 19320 37706 19372
rect 20714 19292 20720 19304
rect 20364 19264 20720 19292
rect 20714 19252 20720 19264
rect 20772 19252 20778 19304
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 21266 19292 21272 19304
rect 20855 19264 21272 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 21266 19252 21272 19264
rect 21324 19252 21330 19304
rect 24210 19292 24216 19304
rect 24171 19264 24216 19292
rect 24210 19252 24216 19264
rect 24268 19252 24274 19304
rect 28350 19292 28356 19304
rect 28311 19264 28356 19292
rect 28350 19252 28356 19264
rect 28408 19252 28414 19304
rect 31386 19292 31392 19304
rect 31347 19264 31392 19292
rect 31386 19252 31392 19264
rect 31444 19252 31450 19304
rect 32493 19295 32551 19301
rect 32493 19261 32505 19295
rect 32539 19292 32551 19295
rect 33226 19292 33232 19304
rect 32539 19264 33232 19292
rect 32539 19261 32551 19264
rect 32493 19255 32551 19261
rect 33226 19252 33232 19264
rect 33284 19252 33290 19304
rect 35526 19292 35532 19304
rect 35487 19264 35532 19292
rect 35526 19252 35532 19264
rect 35584 19252 35590 19304
rect 19702 19156 19708 19168
rect 19663 19128 19708 19156
rect 19702 19116 19708 19128
rect 19760 19116 19766 19168
rect 20717 19159 20775 19165
rect 20717 19125 20729 19159
rect 20763 19156 20775 19159
rect 20806 19156 20812 19168
rect 20763 19128 20812 19156
rect 20763 19125 20775 19128
rect 20717 19119 20775 19125
rect 20806 19116 20812 19128
rect 20864 19156 20870 19168
rect 21634 19156 21640 19168
rect 20864 19128 21640 19156
rect 20864 19116 20870 19128
rect 21634 19116 21640 19128
rect 21692 19116 21698 19168
rect 22370 19116 22376 19168
rect 22428 19156 22434 19168
rect 23385 19159 23443 19165
rect 23385 19156 23397 19159
rect 22428 19128 23397 19156
rect 22428 19116 22434 19128
rect 23385 19125 23397 19128
rect 23431 19125 23443 19159
rect 23385 19119 23443 19125
rect 27157 19159 27215 19165
rect 27157 19125 27169 19159
rect 27203 19156 27215 19159
rect 27246 19156 27252 19168
rect 27203 19128 27252 19156
rect 27203 19125 27215 19128
rect 27157 19119 27215 19125
rect 27246 19116 27252 19128
rect 27304 19116 27310 19168
rect 28445 19159 28503 19165
rect 28445 19125 28457 19159
rect 28491 19156 28503 19159
rect 28718 19156 28724 19168
rect 28491 19128 28724 19156
rect 28491 19125 28503 19128
rect 28445 19119 28503 19125
rect 28718 19116 28724 19128
rect 28776 19116 28782 19168
rect 29273 19159 29331 19165
rect 29273 19125 29285 19159
rect 29319 19156 29331 19159
rect 29822 19156 29828 19168
rect 29319 19128 29828 19156
rect 29319 19125 29331 19128
rect 29273 19119 29331 19125
rect 29822 19116 29828 19128
rect 29880 19116 29886 19168
rect 29914 19116 29920 19168
rect 29972 19156 29978 19168
rect 32490 19156 32496 19168
rect 29972 19128 30017 19156
rect 32451 19128 32496 19156
rect 29972 19116 29978 19128
rect 32490 19116 32496 19128
rect 32548 19116 32554 19168
rect 33318 19116 33324 19168
rect 33376 19156 33382 19168
rect 33413 19159 33471 19165
rect 33413 19156 33425 19159
rect 33376 19128 33425 19156
rect 33376 19116 33382 19128
rect 33413 19125 33425 19128
rect 33459 19125 33471 19159
rect 33413 19119 33471 19125
rect 34517 19159 34575 19165
rect 34517 19125 34529 19159
rect 34563 19156 34575 19159
rect 34698 19156 34704 19168
rect 34563 19128 34704 19156
rect 34563 19125 34575 19128
rect 34517 19119 34575 19125
rect 34698 19116 34704 19128
rect 34756 19116 34762 19168
rect 36630 19116 36636 19168
rect 36688 19156 36694 19168
rect 36909 19159 36967 19165
rect 36909 19156 36921 19159
rect 36688 19128 36921 19156
rect 36688 19116 36694 19128
rect 36909 19125 36921 19128
rect 36955 19125 36967 19159
rect 36909 19119 36967 19125
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 25958 18952 25964 18964
rect 25919 18924 25964 18952
rect 25958 18912 25964 18924
rect 26016 18912 26022 18964
rect 28810 18952 28816 18964
rect 28771 18924 28816 18952
rect 28810 18912 28816 18924
rect 28868 18912 28874 18964
rect 33410 18952 33416 18964
rect 33371 18924 33416 18952
rect 33410 18912 33416 18924
rect 33468 18912 33474 18964
rect 32398 18776 32404 18828
rect 32456 18816 32462 18828
rect 32953 18819 33011 18825
rect 32953 18816 32965 18819
rect 32456 18788 32965 18816
rect 32456 18776 32462 18788
rect 32953 18785 32965 18788
rect 32999 18816 33011 18819
rect 32999 18788 34560 18816
rect 32999 18785 33011 18788
rect 32953 18779 33011 18785
rect 34532 18760 34560 18788
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19613 18751 19671 18757
rect 19613 18748 19625 18751
rect 19484 18720 19625 18748
rect 19484 18708 19490 18720
rect 19613 18717 19625 18720
rect 19659 18717 19671 18751
rect 19613 18711 19671 18717
rect 19702 18708 19708 18760
rect 19760 18748 19766 18760
rect 19869 18751 19927 18757
rect 19869 18748 19881 18751
rect 19760 18720 19881 18748
rect 19760 18708 19766 18720
rect 19869 18717 19881 18720
rect 19915 18717 19927 18751
rect 19869 18711 19927 18717
rect 21266 18708 21272 18760
rect 21324 18748 21330 18760
rect 21453 18751 21511 18757
rect 21453 18748 21465 18751
rect 21324 18720 21465 18748
rect 21324 18708 21330 18720
rect 21453 18717 21465 18720
rect 21499 18717 21511 18751
rect 21634 18748 21640 18760
rect 21595 18720 21640 18748
rect 21453 18711 21511 18717
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 22002 18708 22008 18760
rect 22060 18748 22066 18760
rect 22557 18751 22615 18757
rect 22557 18748 22569 18751
rect 22060 18720 22569 18748
rect 22060 18708 22066 18720
rect 22557 18717 22569 18720
rect 22603 18748 22615 18751
rect 23566 18748 23572 18760
rect 22603 18720 23572 18748
rect 22603 18717 22615 18720
rect 22557 18711 22615 18717
rect 23566 18708 23572 18720
rect 23624 18708 23630 18760
rect 24210 18708 24216 18760
rect 24268 18748 24274 18760
rect 24581 18751 24639 18757
rect 24581 18748 24593 18751
rect 24268 18720 24593 18748
rect 24268 18708 24274 18720
rect 24581 18717 24593 18720
rect 24627 18748 24639 18751
rect 24670 18748 24676 18760
rect 24627 18720 24676 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 24670 18708 24676 18720
rect 24728 18748 24734 18760
rect 26421 18751 26479 18757
rect 26421 18748 26433 18751
rect 24728 18720 26433 18748
rect 24728 18708 24734 18720
rect 26421 18717 26433 18720
rect 26467 18748 26479 18751
rect 27522 18748 27528 18760
rect 26467 18720 27528 18748
rect 26467 18717 26479 18720
rect 26421 18711 26479 18717
rect 27522 18708 27528 18720
rect 27580 18708 27586 18760
rect 28258 18748 28264 18760
rect 28219 18720 28264 18748
rect 28258 18708 28264 18720
rect 28316 18708 28322 18760
rect 28350 18708 28356 18760
rect 28408 18748 28414 18760
rect 28537 18751 28595 18757
rect 28537 18748 28549 18751
rect 28408 18720 28549 18748
rect 28408 18708 28414 18720
rect 28537 18717 28549 18720
rect 28583 18717 28595 18751
rect 31202 18748 31208 18760
rect 31163 18720 31208 18748
rect 28537 18711 28595 18717
rect 31202 18708 31208 18720
rect 31260 18708 31266 18760
rect 33134 18708 33140 18760
rect 33192 18748 33198 18760
rect 33597 18751 33655 18757
rect 33597 18748 33609 18751
rect 33192 18720 33609 18748
rect 33192 18708 33198 18720
rect 33597 18717 33609 18720
rect 33643 18717 33655 18751
rect 34238 18748 34244 18760
rect 34199 18720 34244 18748
rect 33597 18711 33655 18717
rect 34238 18708 34244 18720
rect 34296 18708 34302 18760
rect 34514 18708 34520 18760
rect 34572 18748 34578 18760
rect 34885 18751 34943 18757
rect 34885 18748 34897 18751
rect 34572 18720 34897 18748
rect 34572 18708 34578 18720
rect 34885 18717 34897 18720
rect 34931 18748 34943 18751
rect 35526 18748 35532 18760
rect 34931 18720 35532 18748
rect 34931 18717 34943 18720
rect 34885 18711 34943 18717
rect 35526 18708 35532 18720
rect 35584 18748 35590 18760
rect 36998 18757 37004 18760
rect 36725 18751 36783 18757
rect 36725 18748 36737 18751
rect 35584 18720 36737 18748
rect 35584 18708 35590 18720
rect 36725 18717 36737 18720
rect 36771 18717 36783 18751
rect 36992 18748 37004 18757
rect 36959 18720 37004 18748
rect 36725 18711 36783 18717
rect 36992 18711 37004 18720
rect 36998 18708 37004 18711
rect 37056 18708 37062 18760
rect 19978 18640 19984 18692
rect 20036 18680 20042 18692
rect 20622 18680 20628 18692
rect 20036 18652 20628 18680
rect 20036 18640 20042 18652
rect 20622 18640 20628 18652
rect 20680 18680 20686 18692
rect 21821 18683 21879 18689
rect 21821 18680 21833 18683
rect 20680 18652 21833 18680
rect 20680 18640 20686 18652
rect 21821 18649 21833 18652
rect 21867 18649 21879 18683
rect 21821 18643 21879 18649
rect 22824 18683 22882 18689
rect 22824 18649 22836 18683
rect 22870 18680 22882 18683
rect 23474 18680 23480 18692
rect 22870 18652 23480 18680
rect 22870 18649 22882 18652
rect 22824 18643 22882 18649
rect 23474 18640 23480 18652
rect 23532 18640 23538 18692
rect 24848 18683 24906 18689
rect 24848 18649 24860 18683
rect 24894 18680 24906 18683
rect 25590 18680 25596 18692
rect 24894 18652 25596 18680
rect 24894 18649 24906 18652
rect 24848 18643 24906 18649
rect 25590 18640 25596 18652
rect 25648 18640 25654 18692
rect 26688 18683 26746 18689
rect 26688 18649 26700 18683
rect 26734 18680 26746 18683
rect 28074 18680 28080 18692
rect 26734 18652 28080 18680
rect 26734 18649 26746 18652
rect 26688 18643 26746 18649
rect 28074 18640 28080 18652
rect 28132 18640 28138 18692
rect 28445 18683 28503 18689
rect 28445 18649 28457 18683
rect 28491 18680 28503 18683
rect 28718 18680 28724 18692
rect 28491 18652 28724 18680
rect 28491 18649 28503 18652
rect 28445 18643 28503 18649
rect 28718 18640 28724 18652
rect 28776 18640 28782 18692
rect 34698 18640 34704 18692
rect 34756 18680 34762 18692
rect 35130 18683 35188 18689
rect 35130 18680 35142 18683
rect 34756 18652 35142 18680
rect 34756 18640 34762 18652
rect 35130 18649 35142 18652
rect 35176 18649 35188 18683
rect 35130 18643 35188 18649
rect 20993 18615 21051 18621
rect 20993 18581 21005 18615
rect 21039 18612 21051 18615
rect 21174 18612 21180 18624
rect 21039 18584 21180 18612
rect 21039 18581 21051 18584
rect 20993 18575 21051 18581
rect 21174 18572 21180 18584
rect 21232 18572 21238 18624
rect 23106 18572 23112 18624
rect 23164 18612 23170 18624
rect 23937 18615 23995 18621
rect 23937 18612 23949 18615
rect 23164 18584 23949 18612
rect 23164 18572 23170 18584
rect 23937 18581 23949 18584
rect 23983 18612 23995 18615
rect 25038 18612 25044 18624
rect 23983 18584 25044 18612
rect 23983 18581 23995 18584
rect 23937 18575 23995 18581
rect 25038 18572 25044 18584
rect 25096 18572 25102 18624
rect 27706 18572 27712 18624
rect 27764 18612 27770 18624
rect 27801 18615 27859 18621
rect 27801 18612 27813 18615
rect 27764 18584 27813 18612
rect 27764 18572 27770 18584
rect 27801 18581 27813 18584
rect 27847 18612 27859 18615
rect 28166 18612 28172 18624
rect 27847 18584 28172 18612
rect 27847 18581 27859 18584
rect 27801 18575 27859 18581
rect 28166 18572 28172 18584
rect 28224 18612 28230 18624
rect 28629 18615 28687 18621
rect 28629 18612 28641 18615
rect 28224 18584 28641 18612
rect 28224 18572 28230 18584
rect 28629 18581 28641 18584
rect 28675 18581 28687 18615
rect 34054 18612 34060 18624
rect 34015 18584 34060 18612
rect 28629 18575 28687 18581
rect 34054 18572 34060 18584
rect 34112 18572 34118 18624
rect 36262 18612 36268 18624
rect 36223 18584 36268 18612
rect 36262 18572 36268 18584
rect 36320 18572 36326 18624
rect 37458 18572 37464 18624
rect 37516 18612 37522 18624
rect 38105 18615 38163 18621
rect 38105 18612 38117 18615
rect 37516 18584 38117 18612
rect 37516 18572 37522 18584
rect 38105 18581 38117 18584
rect 38151 18581 38163 18615
rect 38105 18575 38163 18581
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 20162 18408 20168 18420
rect 20123 18380 20168 18408
rect 20162 18368 20168 18380
rect 20220 18368 20226 18420
rect 20806 18368 20812 18420
rect 20864 18417 20870 18420
rect 20864 18411 20883 18417
rect 20871 18377 20883 18411
rect 20864 18371 20883 18377
rect 20864 18368 20870 18371
rect 22186 18368 22192 18420
rect 22244 18408 22250 18420
rect 22649 18411 22707 18417
rect 22649 18408 22661 18411
rect 22244 18380 22661 18408
rect 22244 18368 22250 18380
rect 22649 18377 22661 18380
rect 22695 18377 22707 18411
rect 22649 18371 22707 18377
rect 23566 18368 23572 18420
rect 23624 18408 23630 18420
rect 24673 18411 24731 18417
rect 24673 18408 24685 18411
rect 23624 18380 24685 18408
rect 23624 18368 23630 18380
rect 24673 18377 24685 18380
rect 24719 18377 24731 18411
rect 25590 18408 25596 18420
rect 25551 18380 25596 18408
rect 24673 18371 24731 18377
rect 25590 18368 25596 18380
rect 25648 18368 25654 18420
rect 28350 18368 28356 18420
rect 28408 18408 28414 18420
rect 28537 18411 28595 18417
rect 28537 18408 28549 18411
rect 28408 18380 28549 18408
rect 28408 18368 28414 18380
rect 28537 18377 28549 18380
rect 28583 18377 28595 18411
rect 28537 18371 28595 18377
rect 28810 18368 28816 18420
rect 28868 18408 28874 18420
rect 31113 18411 31171 18417
rect 31113 18408 31125 18411
rect 28868 18380 31125 18408
rect 28868 18368 28874 18380
rect 31113 18377 31125 18380
rect 31159 18377 31171 18411
rect 31113 18371 31171 18377
rect 33226 18368 33232 18420
rect 33284 18408 33290 18420
rect 33781 18411 33839 18417
rect 33781 18408 33793 18411
rect 33284 18380 33793 18408
rect 33284 18368 33290 18380
rect 33781 18377 33793 18380
rect 33827 18377 33839 18411
rect 35986 18408 35992 18420
rect 35947 18380 35992 18408
rect 33781 18371 33839 18377
rect 35986 18368 35992 18380
rect 36044 18368 36050 18420
rect 20625 18343 20683 18349
rect 20625 18340 20637 18343
rect 19904 18312 20637 18340
rect 19904 18281 19932 18312
rect 20625 18309 20637 18312
rect 20671 18340 20683 18343
rect 21174 18340 21180 18352
rect 20671 18312 21180 18340
rect 20671 18309 20683 18312
rect 20625 18303 20683 18309
rect 21174 18300 21180 18312
rect 21232 18300 21238 18352
rect 24118 18340 24124 18352
rect 22664 18312 24124 18340
rect 19889 18275 19947 18281
rect 19889 18241 19901 18275
rect 19935 18241 19947 18275
rect 19889 18235 19947 18241
rect 19978 18232 19984 18284
rect 20036 18272 20042 18284
rect 22370 18272 22376 18284
rect 20036 18244 20081 18272
rect 22331 18244 22376 18272
rect 20036 18232 20042 18244
rect 22370 18232 22376 18244
rect 22428 18232 22434 18284
rect 20165 18207 20223 18213
rect 20165 18173 20177 18207
rect 20211 18204 20223 18207
rect 22094 18204 22100 18216
rect 20211 18176 22100 18204
rect 20211 18173 20223 18176
rect 20165 18167 20223 18173
rect 22094 18164 22100 18176
rect 22152 18204 22158 18216
rect 22664 18213 22692 18312
rect 24118 18300 24124 18312
rect 24176 18300 24182 18352
rect 27522 18340 27528 18352
rect 27172 18312 27528 18340
rect 23382 18272 23388 18284
rect 23295 18244 23388 18272
rect 23382 18232 23388 18244
rect 23440 18232 23446 18284
rect 25774 18272 25780 18284
rect 25735 18244 25780 18272
rect 25774 18232 25780 18244
rect 25832 18232 25838 18284
rect 25958 18232 25964 18284
rect 26016 18272 26022 18284
rect 27172 18281 27200 18312
rect 27522 18300 27528 18312
rect 27580 18300 27586 18352
rect 32668 18343 32726 18349
rect 32668 18309 32680 18343
rect 32714 18340 32726 18343
rect 34054 18340 34060 18352
rect 32714 18312 34060 18340
rect 32714 18309 32726 18312
rect 32668 18303 32726 18309
rect 34054 18300 34060 18312
rect 34112 18300 34118 18352
rect 34698 18340 34704 18352
rect 34659 18312 34704 18340
rect 34698 18300 34704 18312
rect 34756 18300 34762 18352
rect 34793 18343 34851 18349
rect 34793 18309 34805 18343
rect 34839 18340 34851 18343
rect 36262 18340 36268 18352
rect 34839 18312 35480 18340
rect 34839 18309 34851 18312
rect 34793 18303 34851 18309
rect 26053 18275 26111 18281
rect 26053 18272 26065 18275
rect 26016 18244 26065 18272
rect 26016 18232 26022 18244
rect 26053 18241 26065 18244
rect 26099 18241 26111 18275
rect 26053 18235 26111 18241
rect 27157 18275 27215 18281
rect 27157 18241 27169 18275
rect 27203 18241 27215 18275
rect 27157 18235 27215 18241
rect 27246 18232 27252 18284
rect 27304 18272 27310 18284
rect 27413 18275 27471 18281
rect 27413 18272 27425 18275
rect 27304 18244 27425 18272
rect 27304 18232 27310 18244
rect 27413 18241 27425 18244
rect 27459 18241 27471 18275
rect 29730 18272 29736 18284
rect 29691 18244 29736 18272
rect 27413 18235 27471 18241
rect 29730 18232 29736 18244
rect 29788 18232 29794 18284
rect 29822 18232 29828 18284
rect 29880 18272 29886 18284
rect 29989 18275 30047 18281
rect 29989 18272 30001 18275
rect 29880 18244 30001 18272
rect 29880 18232 29886 18244
rect 29989 18241 30001 18244
rect 30035 18241 30047 18275
rect 32398 18272 32404 18284
rect 32359 18244 32404 18272
rect 29989 18235 30047 18241
rect 32398 18232 32404 18244
rect 32456 18232 32462 18284
rect 34609 18275 34667 18281
rect 34609 18241 34621 18275
rect 34655 18241 34667 18275
rect 34911 18275 34969 18281
rect 34911 18272 34923 18275
rect 34609 18235 34667 18241
rect 34716 18244 34923 18272
rect 22649 18207 22707 18213
rect 22649 18204 22661 18207
rect 22152 18176 22661 18204
rect 22152 18164 22158 18176
rect 22649 18173 22661 18176
rect 22695 18173 22707 18207
rect 22649 18167 22707 18173
rect 20714 18096 20720 18148
rect 20772 18136 20778 18148
rect 20993 18139 21051 18145
rect 20993 18136 21005 18139
rect 20772 18108 21005 18136
rect 20772 18096 20778 18108
rect 20993 18105 21005 18108
rect 21039 18105 21051 18139
rect 23400 18136 23428 18232
rect 31202 18136 31208 18148
rect 23400 18108 26096 18136
rect 20993 18099 21051 18105
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 21266 18068 21272 18080
rect 20855 18040 21272 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 21266 18028 21272 18040
rect 21324 18028 21330 18080
rect 22465 18071 22523 18077
rect 22465 18037 22477 18071
rect 22511 18068 22523 18071
rect 24026 18068 24032 18080
rect 22511 18040 24032 18068
rect 22511 18037 22523 18040
rect 22465 18031 22523 18037
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 25130 18028 25136 18080
rect 25188 18068 25194 18080
rect 25866 18068 25872 18080
rect 25188 18040 25872 18068
rect 25188 18028 25194 18040
rect 25866 18028 25872 18040
rect 25924 18068 25930 18080
rect 25961 18071 26019 18077
rect 25961 18068 25973 18071
rect 25924 18040 25973 18068
rect 25924 18028 25930 18040
rect 25961 18037 25973 18040
rect 26007 18037 26019 18071
rect 26068 18068 26096 18108
rect 28092 18108 28672 18136
rect 28092 18068 28120 18108
rect 26068 18040 28120 18068
rect 28644 18068 28672 18108
rect 30668 18108 31208 18136
rect 30668 18068 30696 18108
rect 31202 18096 31208 18108
rect 31260 18096 31266 18148
rect 34624 18136 34652 18235
rect 34716 18216 34744 18244
rect 34911 18241 34923 18244
rect 34957 18241 34969 18275
rect 34911 18235 34969 18241
rect 34698 18164 34704 18216
rect 34756 18164 34762 18216
rect 35069 18207 35127 18213
rect 35069 18173 35081 18207
rect 35115 18204 35127 18207
rect 35342 18204 35348 18216
rect 35115 18176 35348 18204
rect 35115 18173 35127 18176
rect 35069 18167 35127 18173
rect 35342 18164 35348 18176
rect 35400 18164 35406 18216
rect 35452 18204 35480 18312
rect 35728 18312 36268 18340
rect 35728 18281 35756 18312
rect 36262 18300 36268 18312
rect 36320 18340 36326 18352
rect 37461 18343 37519 18349
rect 37461 18340 37473 18343
rect 36320 18312 37473 18340
rect 36320 18300 36326 18312
rect 35713 18275 35771 18281
rect 35713 18241 35725 18275
rect 35759 18241 35771 18275
rect 35713 18235 35771 18241
rect 35805 18275 35863 18281
rect 35805 18241 35817 18275
rect 35851 18272 35863 18275
rect 35894 18272 35900 18284
rect 35851 18244 35900 18272
rect 35851 18241 35863 18244
rect 35805 18235 35863 18241
rect 35894 18232 35900 18244
rect 35952 18232 35958 18284
rect 36648 18281 36676 18312
rect 37461 18309 37473 18312
rect 37507 18309 37519 18343
rect 37461 18303 37519 18309
rect 37550 18300 37556 18352
rect 37608 18340 37614 18352
rect 37661 18343 37719 18349
rect 37661 18340 37673 18343
rect 37608 18312 37673 18340
rect 37608 18300 37614 18312
rect 37661 18309 37673 18312
rect 37707 18309 37719 18343
rect 37661 18303 37719 18309
rect 36449 18275 36507 18281
rect 36449 18241 36461 18275
rect 36495 18241 36507 18275
rect 36449 18235 36507 18241
rect 36633 18275 36691 18281
rect 36633 18241 36645 18275
rect 36679 18241 36691 18275
rect 36633 18235 36691 18241
rect 36464 18204 36492 18235
rect 37458 18204 37464 18216
rect 35452 18176 37464 18204
rect 37458 18164 37464 18176
rect 37516 18164 37522 18216
rect 37829 18139 37887 18145
rect 37829 18136 37841 18139
rect 34624 18108 37841 18136
rect 37829 18105 37841 18108
rect 37875 18105 37887 18139
rect 37829 18099 37887 18105
rect 34422 18068 34428 18080
rect 28644 18040 30696 18068
rect 34383 18040 34428 18068
rect 25961 18031 26019 18037
rect 34422 18028 34428 18040
rect 34480 18028 34486 18080
rect 36538 18068 36544 18080
rect 36499 18040 36544 18068
rect 36538 18028 36544 18040
rect 36596 18028 36602 18080
rect 36814 18068 36820 18080
rect 36775 18040 36820 18068
rect 36814 18028 36820 18040
rect 36872 18028 36878 18080
rect 36906 18028 36912 18080
rect 36964 18068 36970 18080
rect 37645 18071 37703 18077
rect 37645 18068 37657 18071
rect 36964 18040 37657 18068
rect 36964 18028 36970 18040
rect 37645 18037 37657 18040
rect 37691 18037 37703 18071
rect 37645 18031 37703 18037
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 20349 17867 20407 17873
rect 20349 17833 20361 17867
rect 20395 17864 20407 17867
rect 20714 17864 20720 17876
rect 20395 17836 20720 17864
rect 20395 17833 20407 17836
rect 20349 17827 20407 17833
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 22465 17867 22523 17873
rect 22465 17833 22477 17867
rect 22511 17864 22523 17867
rect 23477 17867 23535 17873
rect 22511 17836 22784 17864
rect 22511 17833 22523 17836
rect 22465 17827 22523 17833
rect 20901 17799 20959 17805
rect 20901 17765 20913 17799
rect 20947 17765 20959 17799
rect 20901 17759 20959 17765
rect 20916 17728 20944 17759
rect 21634 17756 21640 17808
rect 21692 17796 21698 17808
rect 22649 17799 22707 17805
rect 22649 17796 22661 17799
rect 21692 17768 22661 17796
rect 21692 17756 21698 17768
rect 22649 17765 22661 17768
rect 22695 17765 22707 17799
rect 22649 17759 22707 17765
rect 20180 17700 20944 17728
rect 20180 17669 20208 17700
rect 20165 17663 20223 17669
rect 20165 17629 20177 17663
rect 20211 17629 20223 17663
rect 20438 17660 20444 17672
rect 20399 17632 20444 17660
rect 20165 17623 20223 17629
rect 20438 17620 20444 17632
rect 20496 17620 20502 17672
rect 20714 17620 20720 17672
rect 20772 17660 20778 17672
rect 21177 17663 21235 17669
rect 21177 17660 21189 17663
rect 20772 17632 21189 17660
rect 20772 17620 20778 17632
rect 21177 17629 21189 17632
rect 21223 17629 21235 17663
rect 21177 17623 21235 17629
rect 22646 17620 22652 17672
rect 22704 17660 22710 17672
rect 22756 17660 22784 17836
rect 23477 17833 23489 17867
rect 23523 17864 23535 17867
rect 24026 17864 24032 17876
rect 23523 17836 24032 17864
rect 23523 17833 23535 17836
rect 23477 17827 23535 17833
rect 24026 17824 24032 17836
rect 24084 17824 24090 17876
rect 25958 17864 25964 17876
rect 25919 17836 25964 17864
rect 25958 17824 25964 17836
rect 26016 17824 26022 17876
rect 26973 17867 27031 17873
rect 26973 17833 26985 17867
rect 27019 17864 27031 17867
rect 27338 17864 27344 17876
rect 27019 17836 27344 17864
rect 27019 17833 27031 17836
rect 26973 17827 27031 17833
rect 27338 17824 27344 17836
rect 27396 17824 27402 17876
rect 28074 17824 28080 17876
rect 28132 17864 28138 17876
rect 29733 17867 29791 17873
rect 29733 17864 29745 17867
rect 28132 17836 29745 17864
rect 28132 17824 28138 17836
rect 29733 17833 29745 17836
rect 29779 17833 29791 17867
rect 29733 17827 29791 17833
rect 29822 17824 29828 17876
rect 29880 17864 29886 17876
rect 32493 17867 32551 17873
rect 32493 17864 32505 17867
rect 29880 17836 32505 17864
rect 29880 17824 29886 17836
rect 32493 17833 32505 17836
rect 32539 17833 32551 17867
rect 32493 17827 32551 17833
rect 33781 17867 33839 17873
rect 33781 17833 33793 17867
rect 33827 17864 33839 17867
rect 34238 17864 34244 17876
rect 33827 17836 34244 17864
rect 33827 17833 33839 17836
rect 33781 17827 33839 17833
rect 34238 17824 34244 17836
rect 34296 17824 34302 17876
rect 35253 17867 35311 17873
rect 35253 17833 35265 17867
rect 35299 17864 35311 17867
rect 35342 17864 35348 17876
rect 35299 17836 35348 17864
rect 35299 17833 35311 17836
rect 35253 17827 35311 17833
rect 35342 17824 35348 17836
rect 35400 17824 35406 17876
rect 36909 17867 36967 17873
rect 36909 17833 36921 17867
rect 36955 17864 36967 17867
rect 37642 17864 37648 17876
rect 36955 17836 37648 17864
rect 36955 17833 36967 17836
rect 36909 17827 36967 17833
rect 37642 17824 37648 17836
rect 37700 17824 37706 17876
rect 25498 17796 25504 17808
rect 24781 17768 25504 17796
rect 23106 17660 23112 17672
rect 22704 17632 23112 17660
rect 22704 17620 22710 17632
rect 23106 17620 23112 17632
rect 23164 17620 23170 17672
rect 23290 17660 23296 17672
rect 23251 17632 23296 17660
rect 23290 17620 23296 17632
rect 23348 17620 23354 17672
rect 24578 17620 24584 17672
rect 24636 17660 24642 17672
rect 24781 17669 24809 17768
rect 25498 17756 25504 17768
rect 25556 17756 25562 17808
rect 28258 17796 28264 17808
rect 27448 17768 28264 17796
rect 27448 17737 27476 17768
rect 28258 17756 28264 17768
rect 28316 17756 28322 17808
rect 35529 17799 35587 17805
rect 35529 17765 35541 17799
rect 35575 17796 35587 17799
rect 36814 17796 36820 17808
rect 35575 17768 36820 17796
rect 35575 17765 35587 17768
rect 35529 17759 35587 17765
rect 36814 17756 36820 17768
rect 36872 17756 36878 17808
rect 26605 17731 26663 17737
rect 25056 17700 25452 17728
rect 24673 17663 24731 17669
rect 24673 17660 24685 17663
rect 24636 17632 24685 17660
rect 24636 17620 24642 17632
rect 24673 17629 24685 17632
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 24766 17663 24824 17669
rect 24766 17629 24778 17663
rect 24812 17629 24824 17663
rect 24766 17623 24824 17629
rect 24903 17663 24961 17669
rect 24903 17629 24915 17663
rect 24949 17660 24961 17663
rect 25056 17660 25084 17700
rect 24949 17632 25084 17660
rect 24949 17629 24961 17632
rect 24903 17623 24961 17629
rect 25130 17620 25136 17672
rect 25188 17669 25194 17672
rect 25188 17660 25196 17669
rect 25188 17632 25233 17660
rect 25188 17623 25196 17632
rect 25188 17620 25194 17623
rect 20898 17592 20904 17604
rect 20859 17564 20904 17592
rect 20898 17552 20904 17564
rect 20956 17552 20962 17604
rect 22186 17552 22192 17604
rect 22244 17592 22250 17604
rect 22281 17595 22339 17601
rect 22281 17592 22293 17595
rect 22244 17564 22293 17592
rect 22244 17552 22250 17564
rect 22281 17561 22293 17564
rect 22327 17592 22339 17595
rect 22370 17592 22376 17604
rect 22327 17564 22376 17592
rect 22327 17561 22339 17564
rect 22281 17555 22339 17561
rect 22370 17552 22376 17564
rect 22428 17552 22434 17604
rect 22497 17595 22555 17601
rect 22497 17561 22509 17595
rect 22543 17592 22555 17595
rect 23308 17592 23336 17620
rect 25424 17604 25452 17700
rect 26605 17697 26617 17731
rect 26651 17697 26663 17731
rect 26605 17691 26663 17697
rect 27433 17731 27491 17737
rect 27433 17697 27445 17731
rect 27479 17697 27491 17731
rect 30377 17731 30435 17737
rect 27433 17691 27491 17697
rect 28644 17700 30052 17728
rect 22543 17564 23336 17592
rect 25041 17595 25099 17601
rect 22543 17561 22555 17564
rect 22497 17555 22555 17561
rect 25041 17561 25053 17595
rect 25087 17592 25099 17595
rect 25222 17592 25228 17604
rect 25087 17564 25228 17592
rect 25087 17561 25099 17564
rect 25041 17555 25099 17561
rect 25222 17552 25228 17564
rect 25280 17552 25286 17604
rect 25406 17552 25412 17604
rect 25464 17592 25470 17604
rect 25777 17595 25835 17601
rect 25777 17592 25789 17595
rect 25464 17564 25789 17592
rect 25464 17552 25470 17564
rect 25777 17561 25789 17564
rect 25823 17561 25835 17595
rect 25777 17555 25835 17561
rect 25866 17552 25872 17604
rect 25924 17592 25930 17604
rect 25977 17595 26035 17601
rect 25977 17592 25989 17595
rect 25924 17564 25989 17592
rect 25924 17552 25930 17564
rect 25977 17561 25989 17564
rect 26023 17592 26035 17595
rect 26510 17592 26516 17604
rect 26023 17564 26516 17592
rect 26023 17561 26035 17564
rect 25977 17555 26035 17561
rect 26510 17552 26516 17564
rect 26568 17552 26574 17604
rect 26620 17592 26648 17691
rect 26786 17660 26792 17672
rect 26747 17632 26792 17660
rect 26786 17620 26792 17632
rect 26844 17660 26850 17672
rect 27617 17663 27675 17669
rect 27617 17660 27629 17663
rect 26844 17632 27629 17660
rect 26844 17620 26850 17632
rect 27617 17629 27629 17632
rect 27663 17660 27675 17663
rect 28644 17660 28672 17700
rect 28810 17660 28816 17672
rect 27663 17632 28672 17660
rect 28771 17632 28816 17660
rect 27663 17629 27675 17632
rect 27617 17623 27675 17629
rect 28810 17620 28816 17632
rect 28868 17620 28874 17672
rect 28920 17669 28948 17700
rect 28905 17663 28963 17669
rect 28905 17629 28917 17663
rect 28951 17629 28963 17663
rect 28905 17623 28963 17629
rect 29917 17663 29975 17669
rect 29917 17629 29929 17663
rect 29963 17629 29975 17663
rect 30024 17660 30052 17700
rect 30377 17697 30389 17731
rect 30423 17728 30435 17731
rect 32490 17728 32496 17740
rect 30423 17700 32496 17728
rect 30423 17697 30435 17700
rect 30377 17691 30435 17697
rect 32490 17688 32496 17700
rect 32548 17688 32554 17740
rect 35452 17700 35894 17728
rect 30558 17660 30564 17672
rect 30024 17632 30564 17660
rect 29917 17623 29975 17629
rect 27706 17592 27712 17604
rect 26620 17564 27712 17592
rect 27706 17552 27712 17564
rect 27764 17552 27770 17604
rect 27801 17595 27859 17601
rect 27801 17561 27813 17595
rect 27847 17592 27859 17595
rect 29932 17592 29960 17623
rect 30558 17620 30564 17632
rect 30616 17620 30622 17672
rect 31202 17660 31208 17672
rect 31163 17632 31208 17660
rect 31202 17620 31208 17632
rect 31260 17620 31266 17672
rect 32306 17620 32312 17672
rect 32364 17660 32370 17672
rect 33410 17660 33416 17672
rect 32364 17632 33416 17660
rect 32364 17620 32370 17632
rect 33410 17620 33416 17632
rect 33468 17620 33474 17672
rect 35452 17669 35480 17700
rect 33597 17663 33655 17669
rect 33597 17629 33609 17663
rect 33643 17629 33655 17663
rect 33597 17623 33655 17629
rect 35437 17663 35495 17669
rect 35437 17629 35449 17663
rect 35483 17629 35495 17663
rect 35437 17623 35495 17629
rect 27847 17564 29960 17592
rect 30576 17592 30604 17620
rect 31570 17592 31576 17604
rect 30576 17564 31576 17592
rect 27847 17561 27859 17564
rect 27801 17555 27859 17561
rect 31570 17552 31576 17564
rect 31628 17592 31634 17604
rect 33612 17592 33640 17623
rect 35526 17620 35532 17672
rect 35584 17660 35590 17672
rect 35621 17663 35679 17669
rect 35621 17660 35633 17663
rect 35584 17632 35633 17660
rect 35584 17620 35590 17632
rect 35621 17629 35633 17632
rect 35667 17629 35679 17663
rect 35749 17663 35807 17669
rect 35749 17660 35761 17663
rect 35621 17623 35679 17629
rect 35728 17629 35761 17660
rect 35795 17629 35807 17663
rect 35866 17660 35894 17700
rect 36630 17660 36636 17672
rect 35866 17632 36636 17660
rect 35728 17623 35807 17629
rect 31628 17564 33640 17592
rect 31628 17552 31634 17564
rect 34790 17552 34796 17604
rect 34848 17592 34854 17604
rect 35728 17592 35756 17623
rect 36630 17620 36636 17632
rect 36688 17620 36694 17672
rect 36725 17663 36783 17669
rect 36725 17629 36737 17663
rect 36771 17629 36783 17663
rect 37458 17660 37464 17672
rect 37419 17632 37464 17660
rect 36725 17623 36783 17629
rect 34848 17564 35756 17592
rect 34848 17552 34854 17564
rect 35894 17552 35900 17604
rect 35952 17592 35958 17604
rect 36740 17592 36768 17623
rect 37458 17620 37464 17632
rect 37516 17620 37522 17672
rect 37553 17663 37611 17669
rect 37553 17629 37565 17663
rect 37599 17629 37611 17663
rect 37553 17623 37611 17629
rect 37568 17592 37596 17623
rect 35952 17564 37596 17592
rect 35952 17552 35958 17564
rect 19978 17524 19984 17536
rect 19939 17496 19984 17524
rect 19978 17484 19984 17496
rect 20036 17484 20042 17536
rect 20438 17484 20444 17536
rect 20496 17524 20502 17536
rect 21085 17527 21143 17533
rect 21085 17524 21097 17527
rect 20496 17496 21097 17524
rect 20496 17484 20502 17496
rect 21085 17493 21097 17496
rect 21131 17493 21143 17527
rect 21085 17487 21143 17493
rect 23658 17484 23664 17536
rect 23716 17524 23722 17536
rect 25317 17527 25375 17533
rect 25317 17524 25329 17527
rect 23716 17496 25329 17524
rect 23716 17484 23722 17496
rect 25317 17493 25329 17496
rect 25363 17493 25375 17527
rect 26142 17524 26148 17536
rect 26103 17496 26148 17524
rect 25317 17487 25375 17493
rect 26142 17484 26148 17496
rect 26200 17484 26206 17536
rect 28994 17484 29000 17536
rect 29052 17524 29058 17536
rect 29089 17527 29147 17533
rect 29089 17524 29101 17527
rect 29052 17496 29101 17524
rect 29052 17484 29058 17496
rect 29089 17493 29101 17496
rect 29135 17493 29147 17527
rect 30742 17524 30748 17536
rect 30703 17496 30748 17524
rect 29089 17487 29147 17493
rect 30742 17484 30748 17496
rect 30800 17484 30806 17536
rect 37642 17484 37648 17536
rect 37700 17524 37706 17536
rect 37737 17527 37795 17533
rect 37737 17524 37749 17527
rect 37700 17496 37749 17524
rect 37700 17484 37706 17496
rect 37737 17493 37749 17496
rect 37783 17493 37795 17527
rect 37737 17487 37795 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 22925 17323 22983 17329
rect 22925 17289 22937 17323
rect 22971 17320 22983 17323
rect 23842 17320 23848 17332
rect 22971 17292 23848 17320
rect 22971 17289 22983 17292
rect 22925 17283 22983 17289
rect 23842 17280 23848 17292
rect 23900 17280 23906 17332
rect 24670 17320 24676 17332
rect 24631 17292 24676 17320
rect 24670 17280 24676 17292
rect 24728 17280 24734 17332
rect 25130 17280 25136 17332
rect 25188 17320 25194 17332
rect 25958 17320 25964 17332
rect 25188 17292 25964 17320
rect 25188 17280 25194 17292
rect 25958 17280 25964 17292
rect 26016 17320 26022 17332
rect 26513 17323 26571 17329
rect 26513 17320 26525 17323
rect 26016 17292 26525 17320
rect 26016 17280 26022 17292
rect 26513 17289 26525 17292
rect 26559 17289 26571 17323
rect 26513 17283 26571 17289
rect 28258 17280 28264 17332
rect 28316 17320 28322 17332
rect 29733 17323 29791 17329
rect 29733 17320 29745 17323
rect 28316 17292 29745 17320
rect 28316 17280 28322 17292
rect 29733 17289 29745 17292
rect 29779 17289 29791 17323
rect 32582 17320 32588 17332
rect 29733 17283 29791 17289
rect 32324 17292 32588 17320
rect 19788 17255 19846 17261
rect 19788 17221 19800 17255
rect 19834 17252 19846 17255
rect 19978 17252 19984 17264
rect 19834 17224 19984 17252
rect 19834 17221 19846 17224
rect 19788 17215 19846 17221
rect 19978 17212 19984 17224
rect 20036 17212 20042 17264
rect 23382 17252 23388 17264
rect 23343 17224 23388 17252
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 25314 17212 25320 17264
rect 25372 17252 25378 17264
rect 26329 17255 26387 17261
rect 26329 17252 26341 17255
rect 25372 17224 26341 17252
rect 25372 17212 25378 17224
rect 26329 17221 26341 17224
rect 26375 17221 26387 17255
rect 27154 17252 27160 17264
rect 27115 17224 27160 17252
rect 26329 17215 26387 17221
rect 27154 17212 27160 17224
rect 27212 17212 27218 17264
rect 27341 17255 27399 17261
rect 27341 17221 27353 17255
rect 27387 17252 27399 17255
rect 27522 17252 27528 17264
rect 27387 17224 27528 17252
rect 27387 17221 27399 17224
rect 27341 17215 27399 17221
rect 27522 17212 27528 17224
rect 27580 17212 27586 17264
rect 28718 17252 28724 17264
rect 28368 17224 28724 17252
rect 19426 17144 19432 17196
rect 19484 17184 19490 17196
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 19484 17156 19533 17184
rect 19484 17144 19490 17156
rect 19521 17153 19533 17156
rect 19567 17153 19579 17187
rect 22646 17184 22652 17196
rect 22607 17156 22652 17184
rect 19521 17147 19579 17153
rect 22646 17144 22652 17156
rect 22704 17144 22710 17196
rect 22741 17187 22799 17193
rect 22741 17153 22753 17187
rect 22787 17184 22799 17187
rect 23290 17184 23296 17196
rect 22787 17156 23296 17184
rect 22787 17153 22799 17156
rect 22741 17147 22799 17153
rect 23290 17144 23296 17156
rect 23348 17184 23354 17196
rect 25593 17187 25651 17193
rect 25593 17184 25605 17187
rect 23348 17156 25605 17184
rect 23348 17144 23354 17156
rect 25593 17153 25605 17156
rect 25639 17184 25651 17187
rect 26142 17184 26148 17196
rect 25639 17156 26148 17184
rect 25639 17153 25651 17156
rect 25593 17147 25651 17153
rect 26142 17144 26148 17156
rect 26200 17144 26206 17196
rect 26510 17144 26516 17196
rect 26568 17184 26574 17196
rect 26605 17187 26663 17193
rect 26605 17184 26617 17187
rect 26568 17156 26617 17184
rect 26568 17144 26574 17156
rect 26605 17153 26617 17156
rect 26651 17153 26663 17187
rect 26605 17147 26663 17153
rect 27246 17144 27252 17196
rect 27304 17184 27310 17196
rect 28368 17193 28396 17224
rect 28718 17212 28724 17224
rect 28776 17252 28782 17264
rect 30466 17261 30472 17264
rect 30460 17252 30472 17261
rect 28776 17224 29776 17252
rect 30427 17224 30472 17252
rect 28776 17212 28782 17224
rect 29748 17196 29776 17224
rect 30460 17215 30472 17224
rect 30466 17212 30472 17215
rect 30524 17212 30530 17264
rect 32214 17212 32220 17264
rect 32272 17252 32278 17264
rect 32324 17261 32352 17292
rect 32582 17280 32588 17292
rect 32640 17280 32646 17332
rect 32858 17320 32864 17332
rect 32819 17292 32864 17320
rect 32858 17280 32864 17292
rect 32916 17280 32922 17332
rect 34790 17320 34796 17332
rect 34751 17292 34796 17320
rect 34790 17280 34796 17292
rect 34848 17280 34854 17332
rect 35526 17280 35532 17332
rect 35584 17320 35590 17332
rect 36817 17323 36875 17329
rect 36817 17320 36829 17323
rect 35584 17292 36829 17320
rect 35584 17280 35590 17292
rect 36817 17289 36829 17292
rect 36863 17289 36875 17323
rect 36817 17283 36875 17289
rect 32309 17255 32367 17261
rect 32309 17252 32321 17255
rect 32272 17224 32321 17252
rect 32272 17212 32278 17224
rect 32309 17221 32321 17224
rect 32355 17221 32367 17255
rect 32490 17252 32496 17264
rect 32451 17224 32496 17252
rect 32309 17215 32367 17221
rect 32490 17212 32496 17224
rect 32548 17212 32554 17264
rect 33226 17252 33232 17264
rect 32600 17224 33232 17252
rect 27433 17187 27491 17193
rect 27433 17184 27445 17187
rect 27304 17156 27445 17184
rect 27304 17144 27310 17156
rect 27433 17153 27445 17156
rect 27479 17153 27491 17187
rect 27433 17147 27491 17153
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17153 28411 17187
rect 28353 17147 28411 17153
rect 28442 17144 28448 17196
rect 28500 17184 28506 17196
rect 28609 17187 28667 17193
rect 28609 17184 28621 17187
rect 28500 17156 28621 17184
rect 28500 17144 28506 17156
rect 28609 17153 28621 17156
rect 28655 17153 28667 17187
rect 28609 17147 28667 17153
rect 29730 17144 29736 17196
rect 29788 17184 29794 17196
rect 30190 17184 30196 17196
rect 29788 17156 30196 17184
rect 29788 17144 29794 17156
rect 30190 17144 30196 17156
rect 30248 17144 30254 17196
rect 32600 17193 32628 17224
rect 33226 17212 33232 17224
rect 33284 17212 33290 17264
rect 33680 17255 33738 17261
rect 33680 17221 33692 17255
rect 33726 17252 33738 17255
rect 34422 17252 34428 17264
rect 33726 17224 34428 17252
rect 33726 17221 33738 17224
rect 33680 17215 33738 17221
rect 34422 17212 34428 17224
rect 34480 17212 34486 17264
rect 36357 17255 36415 17261
rect 36357 17221 36369 17255
rect 36403 17252 36415 17255
rect 37274 17252 37280 17264
rect 36403 17224 37280 17252
rect 36403 17221 36415 17224
rect 36357 17215 36415 17221
rect 37274 17212 37280 17224
rect 37332 17212 37338 17264
rect 32585 17187 32643 17193
rect 32585 17153 32597 17187
rect 32631 17153 32643 17187
rect 32585 17147 32643 17153
rect 32677 17187 32735 17193
rect 32677 17153 32689 17187
rect 32723 17153 32735 17187
rect 35434 17184 35440 17196
rect 35395 17156 35440 17184
rect 32677 17147 32735 17153
rect 22925 17119 22983 17125
rect 22925 17085 22937 17119
rect 22971 17116 22983 17119
rect 24946 17116 24952 17128
rect 22971 17088 24952 17116
rect 22971 17085 22983 17088
rect 22925 17079 22983 17085
rect 24946 17076 24952 17088
rect 25004 17076 25010 17128
rect 25869 17119 25927 17125
rect 25869 17116 25881 17119
rect 25056 17088 25881 17116
rect 24854 17008 24860 17060
rect 24912 17048 24918 17060
rect 25056 17048 25084 17088
rect 25869 17085 25881 17088
rect 25915 17085 25927 17119
rect 25869 17079 25927 17085
rect 32306 17076 32312 17128
rect 32364 17116 32370 17128
rect 32692 17116 32720 17147
rect 35434 17144 35440 17156
rect 35492 17144 35498 17196
rect 36633 17187 36691 17193
rect 36633 17153 36645 17187
rect 36679 17153 36691 17187
rect 37642 17184 37648 17196
rect 37603 17156 37648 17184
rect 36633 17147 36691 17153
rect 32364 17088 32720 17116
rect 33413 17119 33471 17125
rect 32364 17076 32370 17088
rect 33413 17085 33425 17119
rect 33459 17085 33471 17119
rect 33413 17079 33471 17085
rect 24912 17020 25084 17048
rect 25685 17051 25743 17057
rect 24912 17008 24918 17020
rect 25685 17017 25697 17051
rect 25731 17048 25743 17051
rect 26329 17051 26387 17057
rect 26329 17048 26341 17051
rect 25731 17020 26341 17048
rect 25731 17017 25743 17020
rect 25685 17011 25743 17017
rect 26329 17017 26341 17020
rect 26375 17017 26387 17051
rect 26329 17011 26387 17017
rect 31573 17051 31631 17057
rect 31573 17017 31585 17051
rect 31619 17048 31631 17051
rect 32490 17048 32496 17060
rect 31619 17020 32496 17048
rect 31619 17017 31631 17020
rect 31573 17011 31631 17017
rect 32490 17008 32496 17020
rect 32548 17008 32554 17060
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20438 16980 20444 16992
rect 20220 16952 20444 16980
rect 20220 16940 20226 16952
rect 20438 16940 20444 16952
rect 20496 16980 20502 16992
rect 20622 16980 20628 16992
rect 20496 16952 20628 16980
rect 20496 16940 20502 16952
rect 20622 16940 20628 16952
rect 20680 16980 20686 16992
rect 20901 16983 20959 16989
rect 20901 16980 20913 16983
rect 20680 16952 20913 16980
rect 20680 16940 20686 16952
rect 20901 16949 20913 16952
rect 20947 16949 20959 16983
rect 25590 16980 25596 16992
rect 25551 16952 25596 16980
rect 20901 16943 20959 16949
rect 25590 16940 25596 16952
rect 25648 16940 25654 16992
rect 27157 16983 27215 16989
rect 27157 16949 27169 16983
rect 27203 16980 27215 16983
rect 27338 16980 27344 16992
rect 27203 16952 27344 16980
rect 27203 16949 27215 16952
rect 27157 16943 27215 16949
rect 27338 16940 27344 16952
rect 27396 16940 27402 16992
rect 33428 16980 33456 17079
rect 36262 17076 36268 17128
rect 36320 17116 36326 17128
rect 36449 17119 36507 17125
rect 36449 17116 36461 17119
rect 36320 17088 36461 17116
rect 36320 17076 36326 17088
rect 36449 17085 36461 17088
rect 36495 17085 36507 17119
rect 36449 17079 36507 17085
rect 36354 17008 36360 17060
rect 36412 17048 36418 17060
rect 36648 17048 36676 17147
rect 37642 17144 37648 17156
rect 37700 17144 37706 17196
rect 36412 17020 36676 17048
rect 36412 17008 36418 17020
rect 34514 16980 34520 16992
rect 33428 16952 34520 16980
rect 34514 16940 34520 16952
rect 34572 16940 34578 16992
rect 35253 16983 35311 16989
rect 35253 16949 35265 16983
rect 35299 16980 35311 16983
rect 35342 16980 35348 16992
rect 35299 16952 35348 16980
rect 35299 16949 35311 16952
rect 35253 16943 35311 16949
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 36538 16980 36544 16992
rect 36499 16952 36544 16980
rect 36538 16940 36544 16952
rect 36596 16940 36602 16992
rect 37182 16940 37188 16992
rect 37240 16980 37246 16992
rect 37461 16983 37519 16989
rect 37461 16980 37473 16983
rect 37240 16952 37473 16980
rect 37240 16940 37246 16952
rect 37461 16949 37473 16952
rect 37507 16949 37519 16983
rect 37461 16943 37519 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 22186 16736 22192 16788
rect 22244 16776 22250 16788
rect 22244 16748 23612 16776
rect 22244 16736 22250 16748
rect 20438 16668 20444 16720
rect 20496 16668 20502 16720
rect 20622 16668 20628 16720
rect 20680 16668 20686 16720
rect 21266 16668 21272 16720
rect 21324 16708 21330 16720
rect 23474 16708 23480 16720
rect 21324 16680 22094 16708
rect 21324 16668 21330 16680
rect 20456 16640 20484 16668
rect 20456 16612 20576 16640
rect 20254 16572 20260 16584
rect 20215 16544 20260 16572
rect 20254 16532 20260 16544
rect 20312 16532 20318 16584
rect 20548 16581 20576 16612
rect 20640 16581 20668 16668
rect 22066 16640 22094 16680
rect 22480 16680 23480 16708
rect 22373 16643 22431 16649
rect 22373 16640 22385 16643
rect 22066 16612 22385 16640
rect 22373 16609 22385 16612
rect 22419 16609 22431 16643
rect 22373 16603 22431 16609
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16541 20499 16575
rect 20441 16535 20499 16541
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20456 16504 20484 16535
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20809 16575 20867 16581
rect 20809 16572 20821 16575
rect 20772 16544 20821 16572
rect 20772 16532 20778 16544
rect 20809 16541 20821 16544
rect 20855 16541 20867 16575
rect 20809 16535 20867 16541
rect 22005 16575 22063 16581
rect 22005 16541 22017 16575
rect 22051 16541 22063 16575
rect 22186 16572 22192 16584
rect 22147 16544 22192 16572
rect 22005 16535 22063 16541
rect 21174 16504 21180 16516
rect 20456 16476 20668 16504
rect 20640 16436 20668 16476
rect 20824 16476 21180 16504
rect 20824 16436 20852 16476
rect 21174 16464 21180 16476
rect 21232 16464 21238 16516
rect 20990 16436 20996 16448
rect 20640 16408 20852 16436
rect 20951 16408 20996 16436
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 22020 16436 22048 16535
rect 22186 16532 22192 16544
rect 22244 16532 22250 16584
rect 22281 16575 22339 16581
rect 22281 16541 22293 16575
rect 22327 16572 22339 16575
rect 22480 16572 22508 16680
rect 23474 16668 23480 16680
rect 23532 16668 23538 16720
rect 23584 16708 23612 16748
rect 24578 16736 24584 16788
rect 24636 16776 24642 16788
rect 25685 16779 25743 16785
rect 25685 16776 25697 16779
rect 24636 16748 25697 16776
rect 24636 16736 24642 16748
rect 25685 16745 25697 16748
rect 25731 16745 25743 16779
rect 25685 16739 25743 16745
rect 28353 16779 28411 16785
rect 28353 16745 28365 16779
rect 28399 16776 28411 16779
rect 28442 16776 28448 16788
rect 28399 16748 28448 16776
rect 28399 16745 28411 16748
rect 28353 16739 28411 16745
rect 28442 16736 28448 16748
rect 28500 16736 28506 16788
rect 30190 16736 30196 16788
rect 30248 16776 30254 16788
rect 33410 16776 33416 16788
rect 30248 16748 32076 16776
rect 33371 16748 33416 16776
rect 30248 16736 30254 16748
rect 23584 16680 23796 16708
rect 23658 16640 23664 16652
rect 23492 16612 23664 16640
rect 22327 16544 22508 16572
rect 22557 16575 22615 16581
rect 22327 16541 22339 16544
rect 22281 16535 22339 16541
rect 22557 16541 22569 16575
rect 22603 16572 22615 16575
rect 22830 16572 22836 16584
rect 22603 16544 22836 16572
rect 22603 16541 22615 16544
rect 22557 16535 22615 16541
rect 22830 16532 22836 16544
rect 22888 16532 22894 16584
rect 23201 16575 23259 16581
rect 23201 16541 23213 16575
rect 23247 16572 23259 16575
rect 23492 16572 23520 16612
rect 23658 16600 23664 16612
rect 23716 16600 23722 16652
rect 23247 16544 23520 16572
rect 23569 16575 23627 16581
rect 23247 16541 23259 16544
rect 23201 16535 23259 16541
rect 23569 16541 23581 16575
rect 23615 16572 23627 16575
rect 23768 16572 23796 16680
rect 24670 16600 24676 16652
rect 24728 16640 24734 16652
rect 26513 16643 26571 16649
rect 26513 16640 26525 16643
rect 24728 16612 26525 16640
rect 24728 16600 24734 16612
rect 26513 16609 26525 16612
rect 26559 16609 26571 16643
rect 30190 16640 30196 16652
rect 30151 16612 30196 16640
rect 26513 16603 26571 16609
rect 30190 16600 30196 16612
rect 30248 16600 30254 16652
rect 32048 16649 32076 16748
rect 33410 16736 33416 16748
rect 33468 16736 33474 16788
rect 34514 16736 34520 16788
rect 34572 16776 34578 16788
rect 34572 16748 36952 16776
rect 34572 16736 34578 16748
rect 33962 16668 33968 16720
rect 34020 16708 34026 16720
rect 34149 16711 34207 16717
rect 34149 16708 34161 16711
rect 34020 16680 34161 16708
rect 34020 16668 34026 16680
rect 34149 16677 34161 16680
rect 34195 16677 34207 16711
rect 34149 16671 34207 16677
rect 34900 16649 34928 16748
rect 36262 16708 36268 16720
rect 36223 16680 36268 16708
rect 36262 16668 36268 16680
rect 36320 16668 36326 16720
rect 36924 16652 36952 16748
rect 32033 16643 32091 16649
rect 32033 16609 32045 16643
rect 32079 16609 32091 16643
rect 32033 16603 32091 16609
rect 34885 16643 34943 16649
rect 34885 16609 34897 16643
rect 34931 16609 34943 16643
rect 36906 16640 36912 16652
rect 36819 16612 36912 16640
rect 34885 16603 34943 16609
rect 36906 16600 36912 16612
rect 36964 16600 36970 16652
rect 24946 16572 24952 16584
rect 23615 16544 23796 16572
rect 24907 16544 24952 16572
rect 23615 16541 23627 16544
rect 23569 16535 23627 16541
rect 24946 16532 24952 16544
rect 25004 16532 25010 16584
rect 25130 16572 25136 16584
rect 25091 16544 25136 16572
rect 25130 16532 25136 16544
rect 25188 16532 25194 16584
rect 25225 16575 25283 16581
rect 25225 16541 25237 16575
rect 25271 16541 25283 16575
rect 25225 16535 25283 16541
rect 22572 16476 22876 16504
rect 22572 16436 22600 16476
rect 22738 16436 22744 16448
rect 22020 16408 22600 16436
rect 22699 16408 22744 16436
rect 22738 16396 22744 16408
rect 22796 16396 22802 16448
rect 22848 16436 22876 16476
rect 23106 16464 23112 16516
rect 23164 16504 23170 16516
rect 23385 16507 23443 16513
rect 23385 16504 23397 16507
rect 23164 16476 23397 16504
rect 23164 16464 23170 16476
rect 23385 16473 23397 16476
rect 23431 16473 23443 16507
rect 23385 16467 23443 16473
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 25240 16504 25268 16535
rect 25314 16532 25320 16584
rect 25372 16572 25378 16584
rect 25372 16544 25417 16572
rect 25372 16532 25378 16544
rect 25498 16532 25504 16584
rect 25556 16572 25562 16584
rect 28537 16575 28595 16581
rect 25556 16544 25601 16572
rect 25556 16532 25562 16544
rect 28537 16541 28549 16575
rect 28583 16572 28595 16575
rect 28902 16572 28908 16584
rect 28583 16544 28908 16572
rect 28583 16541 28595 16544
rect 28537 16535 28595 16541
rect 28902 16532 28908 16544
rect 28960 16532 28966 16584
rect 28997 16575 29055 16581
rect 28997 16541 29009 16575
rect 29043 16541 29055 16575
rect 28997 16535 29055 16541
rect 33873 16575 33931 16581
rect 33873 16541 33885 16575
rect 33919 16572 33931 16575
rect 34790 16572 34796 16584
rect 33919 16544 34796 16572
rect 33919 16541 33931 16544
rect 33873 16535 33931 16541
rect 25406 16504 25412 16516
rect 23532 16476 23577 16504
rect 25240 16476 25412 16504
rect 23532 16464 23538 16476
rect 25406 16464 25412 16476
rect 25464 16464 25470 16516
rect 26780 16507 26838 16513
rect 26780 16473 26792 16507
rect 26826 16504 26838 16507
rect 27154 16504 27160 16516
rect 26826 16476 27160 16504
rect 26826 16473 26838 16476
rect 26780 16467 26838 16473
rect 27154 16464 27160 16476
rect 27212 16464 27218 16516
rect 29012 16504 29040 16535
rect 34790 16532 34796 16544
rect 34848 16532 34854 16584
rect 37182 16581 37188 16584
rect 37176 16535 37188 16581
rect 37240 16572 37246 16584
rect 37240 16544 37276 16572
rect 37182 16532 37188 16535
rect 37240 16532 37246 16544
rect 27908 16476 29040 16504
rect 30460 16507 30518 16513
rect 23753 16439 23811 16445
rect 23753 16436 23765 16439
rect 22848 16408 23765 16436
rect 23753 16405 23765 16408
rect 23799 16405 23811 16439
rect 23753 16399 23811 16405
rect 27522 16396 27528 16448
rect 27580 16436 27586 16448
rect 27908 16445 27936 16476
rect 30460 16473 30472 16507
rect 30506 16504 30518 16507
rect 30558 16504 30564 16516
rect 30506 16476 30564 16504
rect 30506 16473 30518 16476
rect 30460 16467 30518 16473
rect 30558 16464 30564 16476
rect 30616 16464 30622 16516
rect 30834 16464 30840 16516
rect 30892 16504 30898 16516
rect 32278 16507 32336 16513
rect 32278 16504 32290 16507
rect 30892 16476 32290 16504
rect 30892 16464 30898 16476
rect 32278 16473 32290 16476
rect 32324 16473 32336 16507
rect 32278 16467 32336 16473
rect 35152 16507 35210 16513
rect 35152 16473 35164 16507
rect 35198 16504 35210 16507
rect 35342 16504 35348 16516
rect 35198 16476 35348 16504
rect 35198 16473 35210 16476
rect 35152 16467 35210 16473
rect 35342 16464 35348 16476
rect 35400 16464 35406 16516
rect 27893 16439 27951 16445
rect 27893 16436 27905 16439
rect 27580 16408 27905 16436
rect 27580 16396 27586 16408
rect 27893 16405 27905 16408
rect 27939 16405 27951 16439
rect 29086 16436 29092 16448
rect 29047 16408 29092 16436
rect 27893 16399 27951 16405
rect 29086 16396 29092 16408
rect 29144 16396 29150 16448
rect 31573 16439 31631 16445
rect 31573 16405 31585 16439
rect 31619 16436 31631 16439
rect 32122 16436 32128 16448
rect 31619 16408 32128 16436
rect 31619 16405 31631 16408
rect 31573 16399 31631 16405
rect 32122 16396 32128 16408
rect 32180 16396 32186 16448
rect 34330 16436 34336 16448
rect 34291 16408 34336 16436
rect 34330 16396 34336 16408
rect 34388 16396 34394 16448
rect 37182 16396 37188 16448
rect 37240 16436 37246 16448
rect 38289 16439 38347 16445
rect 38289 16436 38301 16439
rect 37240 16408 38301 16436
rect 37240 16396 37246 16408
rect 38289 16405 38301 16408
rect 38335 16405 38347 16439
rect 38289 16399 38347 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 19705 16235 19763 16241
rect 19705 16201 19717 16235
rect 19751 16232 19763 16235
rect 20622 16232 20628 16244
rect 19751 16204 20628 16232
rect 19751 16201 19763 16204
rect 19705 16195 19763 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 22738 16232 22744 16244
rect 20732 16204 22744 16232
rect 19613 16167 19671 16173
rect 19613 16133 19625 16167
rect 19659 16164 19671 16167
rect 20162 16164 20168 16176
rect 19659 16136 20168 16164
rect 19659 16133 19671 16136
rect 19613 16127 19671 16133
rect 20162 16124 20168 16136
rect 20220 16124 20226 16176
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16096 20039 16099
rect 20070 16096 20076 16108
rect 20027 16068 20076 16096
rect 20027 16065 20039 16068
rect 19981 16059 20039 16065
rect 20070 16056 20076 16068
rect 20128 16056 20134 16108
rect 20732 16105 20760 16204
rect 22738 16192 22744 16204
rect 22796 16192 22802 16244
rect 24946 16192 24952 16244
rect 25004 16232 25010 16244
rect 25501 16235 25559 16241
rect 25501 16232 25513 16235
rect 25004 16204 25513 16232
rect 25004 16192 25010 16204
rect 25501 16201 25513 16204
rect 25547 16201 25559 16235
rect 27154 16232 27160 16244
rect 27115 16204 27160 16232
rect 25501 16195 25559 16201
rect 27154 16192 27160 16204
rect 27212 16192 27218 16244
rect 30558 16232 30564 16244
rect 30519 16204 30564 16232
rect 30558 16192 30564 16204
rect 30616 16192 30622 16244
rect 33226 16232 33232 16244
rect 32968 16204 33232 16232
rect 20993 16167 21051 16173
rect 20993 16133 21005 16167
rect 21039 16164 21051 16167
rect 21266 16164 21272 16176
rect 21039 16136 21272 16164
rect 21039 16133 21051 16136
rect 20993 16127 21051 16133
rect 21266 16124 21272 16136
rect 21324 16124 21330 16176
rect 23928 16167 23986 16173
rect 23928 16133 23940 16167
rect 23974 16164 23986 16167
rect 25590 16164 25596 16176
rect 23974 16136 25596 16164
rect 23974 16133 23986 16136
rect 23928 16127 23986 16133
rect 25590 16124 25596 16136
rect 25648 16124 25654 16176
rect 29086 16164 29092 16176
rect 26068 16136 29092 16164
rect 20898 16105 20904 16108
rect 20717 16099 20775 16105
rect 20717 16065 20729 16099
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 20865 16099 20904 16105
rect 20865 16065 20877 16099
rect 20865 16059 20904 16065
rect 20898 16056 20904 16059
rect 20956 16056 20962 16108
rect 21085 16099 21143 16105
rect 21085 16065 21097 16099
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 20438 15988 20444 16040
rect 20496 16028 20502 16040
rect 21100 16028 21128 16059
rect 21174 16056 21180 16108
rect 21232 16105 21238 16108
rect 21232 16096 21240 16105
rect 21232 16068 21277 16096
rect 21232 16059 21240 16068
rect 21232 16056 21238 16059
rect 22094 16056 22100 16108
rect 22152 16096 22158 16108
rect 22189 16099 22247 16105
rect 22189 16096 22201 16099
rect 22152 16068 22201 16096
rect 22152 16056 22158 16068
rect 22189 16065 22201 16068
rect 22235 16065 22247 16099
rect 22370 16096 22376 16108
rect 22283 16068 22376 16096
rect 22189 16059 22247 16065
rect 22370 16056 22376 16068
rect 22428 16096 22434 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22428 16068 22845 16096
rect 22428 16056 22434 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 23566 16056 23572 16108
rect 23624 16096 23630 16108
rect 23661 16099 23719 16105
rect 23661 16096 23673 16099
rect 23624 16068 23673 16096
rect 23624 16056 23630 16068
rect 23661 16065 23673 16068
rect 23707 16065 23719 16099
rect 23661 16059 23719 16065
rect 25130 16056 25136 16108
rect 25188 16096 25194 16108
rect 25685 16099 25743 16105
rect 25685 16096 25697 16099
rect 25188 16068 25697 16096
rect 25188 16056 25194 16068
rect 25685 16065 25697 16068
rect 25731 16065 25743 16099
rect 25685 16059 25743 16065
rect 25777 16099 25835 16105
rect 25777 16065 25789 16099
rect 25823 16065 25835 16099
rect 25777 16059 25835 16065
rect 25792 16028 25820 16059
rect 25866 16056 25872 16108
rect 25924 16096 25930 16108
rect 26068 16105 26096 16136
rect 29086 16124 29092 16136
rect 29144 16124 29150 16176
rect 25961 16099 26019 16105
rect 25961 16096 25973 16099
rect 25924 16068 25973 16096
rect 25924 16056 25930 16068
rect 25961 16065 25973 16068
rect 26007 16065 26019 16099
rect 25961 16059 26019 16065
rect 26053 16099 26111 16105
rect 26053 16065 26065 16099
rect 26099 16065 26111 16099
rect 27338 16096 27344 16108
rect 27299 16068 27344 16096
rect 26053 16059 26111 16065
rect 27338 16056 27344 16068
rect 27396 16056 27402 16108
rect 27522 16056 27528 16108
rect 27580 16096 27586 16108
rect 27617 16099 27675 16105
rect 27617 16096 27629 16099
rect 27580 16068 27629 16096
rect 27580 16056 27586 16068
rect 27617 16065 27629 16068
rect 27663 16065 27675 16099
rect 27617 16059 27675 16065
rect 28077 16099 28135 16105
rect 28077 16065 28089 16099
rect 28123 16065 28135 16099
rect 28718 16096 28724 16108
rect 28679 16068 28724 16096
rect 28077 16059 28135 16065
rect 20496 16000 21128 16028
rect 25700 16000 25820 16028
rect 28092 16028 28120 16059
rect 28718 16056 28724 16068
rect 28776 16056 28782 16108
rect 28810 16056 28816 16108
rect 28868 16096 28874 16108
rect 28977 16099 29035 16105
rect 28977 16096 28989 16099
rect 28868 16068 28989 16096
rect 28868 16056 28874 16068
rect 28977 16065 28989 16068
rect 29023 16065 29035 16099
rect 30742 16096 30748 16108
rect 30703 16068 30748 16096
rect 28977 16059 29035 16065
rect 30742 16056 30748 16068
rect 30800 16056 30806 16108
rect 31570 16096 31576 16108
rect 31531 16068 31576 16096
rect 31570 16056 31576 16068
rect 31628 16056 31634 16108
rect 32858 16096 32864 16108
rect 32819 16068 32864 16096
rect 32858 16056 32864 16068
rect 32916 16056 32922 16108
rect 32968 16105 32996 16204
rect 33226 16192 33232 16204
rect 33284 16232 33290 16244
rect 34149 16235 34207 16241
rect 34149 16232 34161 16235
rect 33284 16204 34161 16232
rect 33284 16192 33290 16204
rect 34149 16201 34161 16204
rect 34195 16201 34207 16235
rect 34149 16195 34207 16201
rect 35434 16192 35440 16244
rect 35492 16232 35498 16244
rect 35805 16235 35863 16241
rect 35805 16232 35817 16235
rect 35492 16204 35817 16232
rect 35492 16192 35498 16204
rect 35805 16201 35817 16204
rect 35851 16201 35863 16235
rect 35805 16195 35863 16201
rect 36262 16192 36268 16244
rect 36320 16232 36326 16244
rect 36633 16235 36691 16241
rect 36633 16232 36645 16235
rect 36320 16204 36645 16232
rect 36320 16192 36326 16204
rect 36633 16201 36645 16204
rect 36679 16201 36691 16235
rect 36633 16195 36691 16201
rect 36909 16235 36967 16241
rect 36909 16201 36921 16235
rect 36955 16232 36967 16235
rect 37550 16232 37556 16244
rect 36955 16204 37556 16232
rect 36955 16201 36967 16204
rect 36909 16195 36967 16201
rect 37550 16192 37556 16204
rect 37608 16192 37614 16244
rect 36538 16164 36544 16176
rect 36499 16136 36544 16164
rect 36538 16124 36544 16136
rect 36596 16164 36602 16176
rect 37182 16164 37188 16176
rect 36596 16136 37188 16164
rect 36596 16124 36602 16136
rect 37182 16124 37188 16136
rect 37240 16164 37246 16176
rect 37240 16136 37504 16164
rect 37240 16124 37246 16136
rect 32953 16099 33011 16105
rect 32953 16065 32965 16099
rect 32999 16065 33011 16099
rect 32953 16059 33011 16065
rect 33229 16099 33287 16105
rect 33229 16065 33241 16099
rect 33275 16096 33287 16099
rect 33318 16096 33324 16108
rect 33275 16068 33324 16096
rect 33275 16065 33287 16068
rect 33229 16059 33287 16065
rect 33318 16056 33324 16068
rect 33376 16096 33382 16108
rect 34330 16096 34336 16108
rect 33376 16068 34336 16096
rect 33376 16056 33382 16068
rect 34330 16056 34336 16068
rect 34388 16056 34394 16108
rect 35621 16099 35679 16105
rect 35621 16065 35633 16099
rect 35667 16096 35679 16099
rect 35894 16096 35900 16108
rect 35667 16068 35900 16096
rect 35667 16065 35679 16068
rect 35621 16059 35679 16065
rect 35894 16056 35900 16068
rect 35952 16056 35958 16108
rect 36725 16099 36783 16105
rect 36725 16065 36737 16099
rect 36771 16096 36783 16099
rect 37274 16096 37280 16108
rect 36771 16068 37280 16096
rect 36771 16065 36783 16068
rect 36725 16059 36783 16065
rect 31389 16031 31447 16037
rect 28092 16000 28580 16028
rect 20496 15988 20502 16000
rect 19889 15963 19947 15969
rect 19889 15929 19901 15963
rect 19935 15960 19947 15963
rect 20990 15960 20996 15972
rect 19935 15932 20996 15960
rect 19935 15929 19947 15932
rect 19889 15923 19947 15929
rect 20990 15920 20996 15932
rect 21048 15920 21054 15972
rect 21361 15963 21419 15969
rect 21361 15929 21373 15963
rect 21407 15929 21419 15963
rect 21361 15923 21419 15929
rect 25041 15963 25099 15969
rect 25041 15929 25053 15963
rect 25087 15960 25099 15963
rect 25314 15960 25320 15972
rect 25087 15932 25320 15960
rect 25087 15929 25099 15932
rect 25041 15923 25099 15929
rect 19334 15852 19340 15904
rect 19392 15892 19398 15904
rect 19981 15895 20039 15901
rect 19981 15892 19993 15895
rect 19392 15864 19993 15892
rect 19392 15852 19398 15864
rect 19981 15861 19993 15864
rect 20027 15861 20039 15895
rect 19981 15855 20039 15861
rect 20254 15852 20260 15904
rect 20312 15892 20318 15904
rect 21376 15892 21404 15923
rect 25314 15920 25320 15932
rect 25372 15920 25378 15972
rect 25406 15920 25412 15972
rect 25464 15960 25470 15972
rect 25700 15960 25728 16000
rect 28169 15963 28227 15969
rect 28169 15960 28181 15963
rect 25464 15932 28181 15960
rect 25464 15920 25470 15932
rect 28169 15929 28181 15932
rect 28215 15929 28227 15963
rect 28169 15923 28227 15929
rect 20312 15864 21404 15892
rect 22557 15895 22615 15901
rect 20312 15852 20318 15864
rect 22557 15861 22569 15895
rect 22603 15892 22615 15895
rect 26234 15892 26240 15904
rect 22603 15864 26240 15892
rect 22603 15861 22615 15864
rect 22557 15855 22615 15861
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 27525 15895 27583 15901
rect 27525 15861 27537 15895
rect 27571 15892 27583 15895
rect 27890 15892 27896 15904
rect 27571 15864 27896 15892
rect 27571 15861 27583 15864
rect 27525 15855 27583 15861
rect 27890 15852 27896 15864
rect 27948 15852 27954 15904
rect 28552 15892 28580 16000
rect 31389 15997 31401 16031
rect 31435 16028 31447 16031
rect 32122 16028 32128 16040
rect 31435 16000 32128 16028
rect 31435 15997 31447 16000
rect 31389 15991 31447 15997
rect 32122 15988 32128 16000
rect 32180 15988 32186 16040
rect 33689 16031 33747 16037
rect 33689 15997 33701 16031
rect 33735 16028 33747 16031
rect 33962 16028 33968 16040
rect 33735 16000 33968 16028
rect 33735 15997 33747 16000
rect 33689 15991 33747 15997
rect 31478 15920 31484 15972
rect 31536 15960 31542 15972
rect 33704 15960 33732 15991
rect 33962 15988 33968 16000
rect 34020 15988 34026 16040
rect 35437 16031 35495 16037
rect 35437 15997 35449 16031
rect 35483 16028 35495 16031
rect 36740 16028 36768 16059
rect 37274 16056 37280 16068
rect 37332 16056 37338 16108
rect 37476 16105 37504 16136
rect 37461 16099 37519 16105
rect 37461 16065 37473 16099
rect 37507 16065 37519 16099
rect 37642 16096 37648 16108
rect 37603 16068 37648 16096
rect 37461 16059 37519 16065
rect 37642 16056 37648 16068
rect 37700 16056 37706 16108
rect 35483 16000 36768 16028
rect 35483 15997 35495 16000
rect 35437 15991 35495 15997
rect 31536 15932 33732 15960
rect 34057 15963 34115 15969
rect 31536 15920 31542 15932
rect 34057 15929 34069 15963
rect 34103 15960 34115 15963
rect 34790 15960 34796 15972
rect 34103 15932 34796 15960
rect 34103 15929 34115 15932
rect 34057 15923 34115 15929
rect 34790 15920 34796 15932
rect 34848 15920 34854 15972
rect 36170 15920 36176 15972
rect 36228 15960 36234 15972
rect 36354 15960 36360 15972
rect 36228 15932 36360 15960
rect 36228 15920 36234 15932
rect 36354 15920 36360 15932
rect 36412 15920 36418 15972
rect 29362 15892 29368 15904
rect 28552 15864 29368 15892
rect 29362 15852 29368 15864
rect 29420 15892 29426 15904
rect 30101 15895 30159 15901
rect 30101 15892 30113 15895
rect 29420 15864 30113 15892
rect 29420 15852 29426 15864
rect 30101 15861 30113 15864
rect 30147 15861 30159 15895
rect 30101 15855 30159 15861
rect 30926 15852 30932 15904
rect 30984 15892 30990 15904
rect 31757 15895 31815 15901
rect 31757 15892 31769 15895
rect 30984 15864 31769 15892
rect 30984 15852 30990 15864
rect 31757 15861 31769 15864
rect 31803 15861 31815 15895
rect 32674 15892 32680 15904
rect 32635 15864 32680 15892
rect 31757 15855 31815 15861
rect 32674 15852 32680 15864
rect 32732 15852 32738 15904
rect 33134 15892 33140 15904
rect 33095 15864 33140 15892
rect 33134 15852 33140 15864
rect 33192 15852 33198 15904
rect 37829 15895 37887 15901
rect 37829 15861 37841 15895
rect 37875 15892 37887 15895
rect 38286 15892 38292 15904
rect 37875 15864 38292 15892
rect 37875 15861 37887 15864
rect 37829 15855 37887 15861
rect 38286 15852 38292 15864
rect 38344 15852 38350 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1854 15648 1860 15700
rect 1912 15688 1918 15700
rect 20438 15688 20444 15700
rect 1912 15660 6914 15688
rect 20399 15660 20444 15688
rect 1912 15648 1918 15660
rect 6886 15620 6914 15660
rect 20438 15648 20444 15660
rect 20496 15648 20502 15700
rect 20898 15648 20904 15700
rect 20956 15688 20962 15700
rect 22189 15691 22247 15697
rect 22189 15688 22201 15691
rect 20956 15660 22201 15688
rect 20956 15648 20962 15660
rect 22189 15657 22201 15660
rect 22235 15688 22247 15691
rect 22830 15688 22836 15700
rect 22235 15660 22836 15688
rect 22235 15657 22247 15660
rect 22189 15651 22247 15657
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 23106 15688 23112 15700
rect 23067 15660 23112 15688
rect 23106 15648 23112 15660
rect 23164 15648 23170 15700
rect 23474 15648 23480 15700
rect 23532 15688 23538 15700
rect 23661 15691 23719 15697
rect 23661 15688 23673 15691
rect 23532 15660 23673 15688
rect 23532 15648 23538 15660
rect 23661 15657 23673 15660
rect 23707 15657 23719 15691
rect 23661 15651 23719 15657
rect 26789 15691 26847 15697
rect 26789 15657 26801 15691
rect 26835 15688 26847 15691
rect 27798 15688 27804 15700
rect 26835 15660 27804 15688
rect 26835 15657 26847 15660
rect 26789 15651 26847 15657
rect 27798 15648 27804 15660
rect 27856 15648 27862 15700
rect 28445 15691 28503 15697
rect 28445 15657 28457 15691
rect 28491 15688 28503 15691
rect 28810 15688 28816 15700
rect 28491 15660 28816 15688
rect 28491 15657 28503 15660
rect 28445 15651 28503 15657
rect 28810 15648 28816 15660
rect 28868 15648 28874 15700
rect 29086 15648 29092 15700
rect 29144 15688 29150 15700
rect 30374 15688 30380 15700
rect 29144 15660 30380 15688
rect 29144 15648 29150 15660
rect 30374 15648 30380 15660
rect 30432 15648 30438 15700
rect 30745 15691 30803 15697
rect 30745 15657 30757 15691
rect 30791 15688 30803 15691
rect 30834 15688 30840 15700
rect 30791 15660 30840 15688
rect 30791 15657 30803 15660
rect 30745 15651 30803 15657
rect 30834 15648 30840 15660
rect 30892 15648 30898 15700
rect 33226 15688 33232 15700
rect 33187 15660 33232 15688
rect 33226 15648 33232 15660
rect 33284 15648 33290 15700
rect 36170 15648 36176 15700
rect 36228 15688 36234 15700
rect 38289 15691 38347 15697
rect 38289 15688 38301 15691
rect 36228 15660 38301 15688
rect 36228 15648 36234 15660
rect 38289 15657 38301 15660
rect 38335 15657 38347 15691
rect 38289 15651 38347 15657
rect 22370 15620 22376 15632
rect 6886 15592 22376 15620
rect 22370 15580 22376 15592
rect 22428 15580 22434 15632
rect 27433 15623 27491 15629
rect 27433 15620 27445 15623
rect 26712 15592 27445 15620
rect 20349 15487 20407 15493
rect 20349 15453 20361 15487
rect 20395 15453 20407 15487
rect 20349 15447 20407 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15484 21051 15487
rect 21174 15484 21180 15496
rect 21039 15456 21180 15484
rect 21039 15453 21051 15456
rect 20993 15447 21051 15453
rect 20364 15416 20392 15447
rect 21174 15444 21180 15456
rect 21232 15444 21238 15496
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22152 15456 22197 15484
rect 22152 15444 22158 15456
rect 22646 15444 22652 15496
rect 22704 15484 22710 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22704 15456 22753 15484
rect 22704 15444 22710 15456
rect 22741 15453 22753 15456
rect 22787 15453 22799 15487
rect 22741 15447 22799 15453
rect 23569 15487 23627 15493
rect 23569 15453 23581 15487
rect 23615 15484 23627 15487
rect 23658 15484 23664 15496
rect 23615 15456 23664 15484
rect 23615 15453 23627 15456
rect 23569 15447 23627 15453
rect 23658 15444 23664 15456
rect 23716 15484 23722 15496
rect 25314 15484 25320 15496
rect 23716 15456 25320 15484
rect 23716 15444 23722 15456
rect 25314 15444 25320 15456
rect 25372 15444 25378 15496
rect 26712 15493 26740 15592
rect 27433 15589 27445 15592
rect 27479 15589 27491 15623
rect 35894 15620 35900 15632
rect 27433 15583 27491 15589
rect 27540 15592 29224 15620
rect 26973 15555 27031 15561
rect 26973 15521 26985 15555
rect 27019 15552 27031 15555
rect 27246 15552 27252 15564
rect 27019 15524 27252 15552
rect 27019 15521 27031 15524
rect 26973 15515 27031 15521
rect 27246 15512 27252 15524
rect 27304 15552 27310 15564
rect 27540 15552 27568 15592
rect 27304 15524 27568 15552
rect 27304 15512 27310 15524
rect 27890 15512 27896 15564
rect 27948 15552 27954 15564
rect 27948 15524 28856 15552
rect 27948 15512 27954 15524
rect 26697 15487 26755 15493
rect 26697 15453 26709 15487
rect 26743 15453 26755 15487
rect 26697 15447 26755 15453
rect 26988 15456 27660 15484
rect 21450 15416 21456 15428
rect 20364 15388 21456 15416
rect 21450 15376 21456 15388
rect 21508 15376 21514 15428
rect 22925 15419 22983 15425
rect 22925 15385 22937 15419
rect 22971 15416 22983 15419
rect 25222 15416 25228 15428
rect 22971 15388 25228 15416
rect 22971 15385 22983 15388
rect 22925 15379 22983 15385
rect 25222 15376 25228 15388
rect 25280 15416 25286 15428
rect 25866 15416 25872 15428
rect 25280 15388 25872 15416
rect 25280 15376 25286 15388
rect 25866 15376 25872 15388
rect 25924 15376 25930 15428
rect 26988 15425 27016 15456
rect 26973 15419 27031 15425
rect 26973 15385 26985 15419
rect 27019 15385 27031 15419
rect 26973 15379 27031 15385
rect 27433 15419 27491 15425
rect 27433 15385 27445 15419
rect 27479 15416 27491 15419
rect 27522 15416 27528 15428
rect 27479 15388 27528 15416
rect 27479 15385 27491 15388
rect 27433 15379 27491 15385
rect 27522 15376 27528 15388
rect 27580 15376 27586 15428
rect 27632 15416 27660 15456
rect 27706 15444 27712 15496
rect 27764 15484 27770 15496
rect 27764 15456 27809 15484
rect 27764 15444 27770 15456
rect 28534 15444 28540 15496
rect 28592 15486 28598 15496
rect 28828 15493 28856 15524
rect 28701 15487 28759 15493
rect 28701 15486 28713 15487
rect 28592 15458 28713 15486
rect 28592 15444 28598 15458
rect 28701 15453 28713 15458
rect 28747 15453 28759 15487
rect 28701 15447 28759 15453
rect 28813 15487 28871 15493
rect 28813 15453 28825 15487
rect 28859 15453 28871 15487
rect 28813 15447 28871 15453
rect 28905 15487 28963 15493
rect 28905 15453 28917 15487
rect 28951 15453 28963 15487
rect 29086 15484 29092 15496
rect 29047 15456 29092 15484
rect 28905 15447 28963 15453
rect 28933 15416 28961 15447
rect 29086 15444 29092 15456
rect 29144 15444 29150 15496
rect 27632 15388 28961 15416
rect 29196 15416 29224 15592
rect 35866 15580 35900 15620
rect 35952 15620 35958 15632
rect 35952 15592 36308 15620
rect 35952 15580 35958 15592
rect 31757 15555 31815 15561
rect 31757 15552 31769 15555
rect 30300 15524 31769 15552
rect 30300 15493 30328 15524
rect 31757 15521 31769 15524
rect 31803 15521 31815 15555
rect 33134 15552 33140 15564
rect 31757 15515 31815 15521
rect 32968 15524 33140 15552
rect 30285 15487 30343 15493
rect 30285 15453 30297 15487
rect 30331 15453 30343 15487
rect 30926 15484 30932 15496
rect 30887 15456 30932 15484
rect 30285 15447 30343 15453
rect 30926 15444 30932 15456
rect 30984 15444 30990 15496
rect 31478 15484 31484 15496
rect 31439 15456 31484 15484
rect 31478 15444 31484 15456
rect 31536 15444 31542 15496
rect 32968 15493 32996 15524
rect 33134 15512 33140 15524
rect 33192 15512 33198 15564
rect 33318 15552 33324 15564
rect 33279 15524 33324 15552
rect 33318 15512 33324 15524
rect 33376 15512 33382 15564
rect 33781 15555 33839 15561
rect 33781 15521 33793 15555
rect 33827 15552 33839 15555
rect 34790 15552 34796 15564
rect 33827 15524 34796 15552
rect 33827 15521 33839 15524
rect 33781 15515 33839 15521
rect 34790 15512 34796 15524
rect 34848 15512 34854 15564
rect 31573 15487 31631 15493
rect 31573 15453 31585 15487
rect 31619 15484 31631 15487
rect 32953 15487 33011 15493
rect 31619 15456 31754 15484
rect 31619 15453 31631 15456
rect 31573 15447 31631 15453
rect 31726 15416 31754 15456
rect 32953 15453 32965 15487
rect 32999 15453 33011 15487
rect 32953 15447 33011 15453
rect 33042 15444 33048 15496
rect 33100 15484 33106 15496
rect 33965 15487 34023 15493
rect 33100 15456 33145 15484
rect 33100 15444 33106 15456
rect 33965 15453 33977 15487
rect 34011 15453 34023 15487
rect 33965 15447 34023 15453
rect 34149 15487 34207 15493
rect 34149 15453 34161 15487
rect 34195 15484 34207 15487
rect 35069 15487 35127 15493
rect 35069 15484 35081 15487
rect 34195 15456 35081 15484
rect 34195 15453 34207 15456
rect 34149 15447 34207 15453
rect 35069 15453 35081 15456
rect 35115 15453 35127 15487
rect 35069 15447 35127 15453
rect 33980 15416 34008 15447
rect 35866 15416 35894 15580
rect 36170 15484 36176 15496
rect 36131 15456 36176 15484
rect 36170 15444 36176 15456
rect 36228 15444 36234 15496
rect 36280 15493 36308 15592
rect 36906 15552 36912 15564
rect 36867 15524 36912 15552
rect 36906 15512 36912 15524
rect 36964 15512 36970 15564
rect 36265 15487 36323 15493
rect 36265 15453 36277 15487
rect 36311 15484 36323 15487
rect 37642 15484 37648 15496
rect 36311 15456 37648 15484
rect 36311 15453 36323 15456
rect 36265 15447 36323 15453
rect 37642 15444 37648 15456
rect 37700 15444 37706 15496
rect 29196 15388 30788 15416
rect 31726 15388 35894 15416
rect 37176 15419 37234 15425
rect 21177 15351 21235 15357
rect 21177 15317 21189 15351
rect 21223 15348 21235 15351
rect 21358 15348 21364 15360
rect 21223 15320 21364 15348
rect 21223 15317 21235 15320
rect 21177 15311 21235 15317
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 27614 15348 27620 15360
rect 27575 15320 27620 15348
rect 27614 15308 27620 15320
rect 27672 15308 27678 15360
rect 28902 15308 28908 15360
rect 28960 15348 28966 15360
rect 29362 15348 29368 15360
rect 28960 15320 29368 15348
rect 28960 15308 28966 15320
rect 29362 15308 29368 15320
rect 29420 15308 29426 15360
rect 30101 15351 30159 15357
rect 30101 15317 30113 15351
rect 30147 15348 30159 15351
rect 30650 15348 30656 15360
rect 30147 15320 30656 15348
rect 30147 15317 30159 15320
rect 30101 15311 30159 15317
rect 30650 15308 30656 15320
rect 30708 15308 30714 15360
rect 30760 15348 30788 15388
rect 37176 15385 37188 15419
rect 37222 15416 37234 15419
rect 38102 15416 38108 15428
rect 37222 15388 38108 15416
rect 37222 15385 37234 15388
rect 37176 15379 37234 15385
rect 38102 15376 38108 15388
rect 38160 15376 38166 15428
rect 32769 15351 32827 15357
rect 32769 15348 32781 15351
rect 30760 15320 32781 15348
rect 32769 15317 32781 15320
rect 32815 15317 32827 15351
rect 34882 15348 34888 15360
rect 34843 15320 34888 15348
rect 32769 15311 32827 15317
rect 34882 15308 34888 15320
rect 34940 15308 34946 15360
rect 36449 15351 36507 15357
rect 36449 15317 36461 15351
rect 36495 15348 36507 15351
rect 37642 15348 37648 15360
rect 36495 15320 37648 15348
rect 36495 15317 36507 15320
rect 36449 15311 36507 15317
rect 37642 15308 37648 15320
rect 37700 15308 37706 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22738 15144 22744 15156
rect 22152 15116 22744 15144
rect 22152 15104 22158 15116
rect 22738 15104 22744 15116
rect 22796 15144 22802 15156
rect 23477 15147 23535 15153
rect 23477 15144 23489 15147
rect 22796 15116 23489 15144
rect 22796 15104 22802 15116
rect 23477 15113 23489 15116
rect 23523 15113 23535 15147
rect 25314 15144 25320 15156
rect 25275 15116 25320 15144
rect 23477 15107 23535 15113
rect 25314 15104 25320 15116
rect 25372 15104 25378 15156
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 26513 15147 26571 15153
rect 26513 15144 26525 15147
rect 25556 15116 26525 15144
rect 25556 15104 25562 15116
rect 26513 15113 26525 15116
rect 26559 15113 26571 15147
rect 27706 15144 27712 15156
rect 26513 15107 26571 15113
rect 27172 15116 27712 15144
rect 23566 15076 23572 15088
rect 20088 15048 23572 15076
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 20088 15017 20116 15048
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19484 14980 20085 15008
rect 19484 14968 19490 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20340 15011 20398 15017
rect 20340 14977 20352 15011
rect 20386 15008 20398 15011
rect 21266 15008 21272 15020
rect 20386 14980 21272 15008
rect 20386 14977 20398 14980
rect 20340 14971 20398 14977
rect 21266 14968 21272 14980
rect 21324 14968 21330 15020
rect 22112 15017 22140 15048
rect 23566 15036 23572 15048
rect 23624 15036 23630 15088
rect 24670 15076 24676 15088
rect 23952 15048 24676 15076
rect 22097 15011 22155 15017
rect 22097 14977 22109 15011
rect 22143 15008 22155 15011
rect 22364 15011 22422 15017
rect 22143 14980 22177 15008
rect 22143 14977 22155 14980
rect 22097 14971 22155 14977
rect 22364 14977 22376 15011
rect 22410 15008 22422 15011
rect 22922 15008 22928 15020
rect 22410 14980 22928 15008
rect 22410 14977 22422 14980
rect 22364 14971 22422 14977
rect 22922 14968 22928 14980
rect 22980 14968 22986 15020
rect 23952 15017 23980 15048
rect 24670 15036 24676 15048
rect 24728 15036 24734 15088
rect 25866 15076 25872 15088
rect 25827 15048 25872 15076
rect 25866 15036 25872 15048
rect 25924 15036 25930 15088
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 24026 14968 24032 15020
rect 24084 15008 24090 15020
rect 24193 15011 24251 15017
rect 24193 15008 24205 15011
rect 24084 14980 24205 15008
rect 24084 14968 24090 14980
rect 24193 14977 24205 14980
rect 24239 14977 24251 15011
rect 24193 14971 24251 14977
rect 25777 15011 25835 15017
rect 25777 14977 25789 15011
rect 25823 15008 25835 15011
rect 26326 15008 26332 15020
rect 25823 14980 26332 15008
rect 25823 14977 25835 14980
rect 25777 14971 25835 14977
rect 26326 14968 26332 14980
rect 26384 14968 26390 15020
rect 26418 14968 26424 15020
rect 26476 15008 26482 15020
rect 27172 15017 27200 15116
rect 27706 15104 27712 15116
rect 27764 15144 27770 15156
rect 28997 15147 29055 15153
rect 28997 15144 29009 15147
rect 27764 15116 29009 15144
rect 27764 15104 27770 15116
rect 28997 15113 29009 15116
rect 29043 15113 29055 15147
rect 28997 15107 29055 15113
rect 31386 15104 31392 15156
rect 31444 15144 31450 15156
rect 31573 15147 31631 15153
rect 31573 15144 31585 15147
rect 31444 15116 31585 15144
rect 31444 15104 31450 15116
rect 31573 15113 31585 15116
rect 31619 15113 31631 15147
rect 33134 15144 33140 15156
rect 33095 15116 33140 15144
rect 31573 15107 31631 15113
rect 33134 15104 33140 15116
rect 33192 15104 33198 15156
rect 34977 15147 35035 15153
rect 34977 15144 34989 15147
rect 33520 15116 34989 15144
rect 27522 15076 27528 15088
rect 27483 15048 27528 15076
rect 27522 15036 27528 15048
rect 27580 15036 27586 15088
rect 28445 15079 28503 15085
rect 28445 15076 28457 15079
rect 27632 15048 28457 15076
rect 27632 15020 27660 15048
rect 28445 15045 28457 15048
rect 28491 15045 28503 15079
rect 28445 15039 28503 15045
rect 28624 15048 29132 15076
rect 27157 15011 27215 15017
rect 26476 14980 26521 15008
rect 26476 14968 26482 14980
rect 27157 14977 27169 15011
rect 27203 14977 27215 15011
rect 27157 14971 27215 14977
rect 27614 14968 27620 15020
rect 27672 15008 27678 15020
rect 28077 15011 28135 15017
rect 27672 14980 27765 15008
rect 27672 14968 27678 14980
rect 28077 14977 28089 15011
rect 28123 14977 28135 15011
rect 28077 14971 28135 14977
rect 28261 15011 28319 15017
rect 28261 14977 28273 15011
rect 28307 15008 28319 15011
rect 28624 15008 28652 15048
rect 28902 15008 28908 15020
rect 28307 14980 28652 15008
rect 28863 14980 28908 15008
rect 28307 14977 28319 14980
rect 28261 14971 28319 14977
rect 28092 14884 28120 14971
rect 28902 14968 28908 14980
rect 28960 14968 28966 15020
rect 29104 15017 29132 15048
rect 29089 15011 29147 15017
rect 29089 14977 29101 15011
rect 29135 15008 29147 15011
rect 29362 15008 29368 15020
rect 29135 14980 29368 15008
rect 29135 14977 29147 14980
rect 29089 14971 29147 14977
rect 29362 14968 29368 14980
rect 29420 14968 29426 15020
rect 30006 14968 30012 15020
rect 30064 15008 30070 15020
rect 30449 15011 30507 15017
rect 30449 15008 30461 15011
rect 30064 14980 30461 15008
rect 30064 14968 30070 14980
rect 30449 14977 30461 14980
rect 30495 14977 30507 15011
rect 30449 14971 30507 14977
rect 32953 15011 33011 15017
rect 32953 14977 32965 15011
rect 32999 15008 33011 15011
rect 33042 15008 33048 15020
rect 32999 14980 33048 15008
rect 32999 14977 33011 14980
rect 32953 14971 33011 14977
rect 33042 14968 33048 14980
rect 33100 15008 33106 15020
rect 33520 15008 33548 15116
rect 34977 15113 34989 15116
rect 35023 15113 35035 15147
rect 34977 15107 35035 15113
rect 36630 15104 36636 15156
rect 36688 15144 36694 15156
rect 36817 15147 36875 15153
rect 36817 15144 36829 15147
rect 36688 15116 36829 15144
rect 36688 15104 36694 15116
rect 36817 15113 36829 15116
rect 36863 15113 36875 15147
rect 38102 15144 38108 15156
rect 38063 15116 38108 15144
rect 36817 15107 36875 15113
rect 38102 15104 38108 15116
rect 38160 15104 38166 15156
rect 35894 15076 35900 15088
rect 33612 15048 35900 15076
rect 33612 15017 33640 15048
rect 33100 14980 33548 15008
rect 33597 15011 33655 15017
rect 33100 14968 33106 14980
rect 33597 14977 33609 15011
rect 33643 14977 33655 15011
rect 33597 14971 33655 14977
rect 33864 15011 33922 15017
rect 33864 14977 33876 15011
rect 33910 15008 33922 15011
rect 34882 15008 34888 15020
rect 33910 14980 34888 15008
rect 33910 14977 33922 14980
rect 33864 14971 33922 14977
rect 34882 14968 34888 14980
rect 34940 14968 34946 15020
rect 35452 15017 35480 15048
rect 35894 15036 35900 15048
rect 35952 15076 35958 15088
rect 36906 15076 36912 15088
rect 35952 15048 36912 15076
rect 35952 15036 35958 15048
rect 36906 15036 36912 15048
rect 36964 15036 36970 15088
rect 35437 15011 35495 15017
rect 35437 14977 35449 15011
rect 35483 14977 35495 15011
rect 35437 14971 35495 14977
rect 35526 14968 35532 15020
rect 35584 15008 35590 15020
rect 35693 15011 35751 15017
rect 35693 15008 35705 15011
rect 35584 14980 35705 15008
rect 35584 14968 35590 14980
rect 35693 14977 35705 14980
rect 35739 14977 35751 15011
rect 37642 15008 37648 15020
rect 37603 14980 37648 15008
rect 35693 14971 35751 14977
rect 37642 14968 37648 14980
rect 37700 14968 37706 15020
rect 38286 15008 38292 15020
rect 38247 14980 38292 15008
rect 38286 14968 38292 14980
rect 38344 14968 38350 15020
rect 28718 14900 28724 14952
rect 28776 14940 28782 14952
rect 30193 14943 30251 14949
rect 30193 14940 30205 14943
rect 28776 14912 30205 14940
rect 28776 14900 28782 14912
rect 30193 14909 30205 14912
rect 30239 14909 30251 14943
rect 30193 14903 30251 14909
rect 32582 14900 32588 14952
rect 32640 14940 32646 14952
rect 32769 14943 32827 14949
rect 32769 14940 32781 14943
rect 32640 14912 32781 14940
rect 32640 14900 32646 14912
rect 32769 14909 32781 14912
rect 32815 14909 32827 14943
rect 32769 14903 32827 14909
rect 28074 14872 28080 14884
rect 27987 14844 28080 14872
rect 28074 14832 28080 14844
rect 28132 14872 28138 14884
rect 28132 14844 28948 14872
rect 28132 14832 28138 14844
rect 28920 14816 28948 14844
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 27338 14804 27344 14816
rect 27299 14776 27344 14804
rect 27338 14764 27344 14776
rect 27396 14764 27402 14816
rect 28902 14764 28908 14816
rect 28960 14804 28966 14816
rect 32674 14804 32680 14816
rect 28960 14776 32680 14804
rect 28960 14764 28966 14776
rect 32674 14764 32680 14776
rect 32732 14764 32738 14816
rect 37458 14804 37464 14816
rect 37419 14776 37464 14804
rect 37458 14764 37464 14776
rect 37516 14764 37522 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 21266 14600 21272 14612
rect 21227 14572 21272 14600
rect 21266 14560 21272 14572
rect 21324 14560 21330 14612
rect 23385 14603 23443 14609
rect 23385 14569 23397 14603
rect 23431 14600 23443 14603
rect 24026 14600 24032 14612
rect 23431 14572 24032 14600
rect 23431 14569 23443 14572
rect 23385 14563 23443 14569
rect 24026 14560 24032 14572
rect 24084 14560 24090 14612
rect 27614 14600 27620 14612
rect 27575 14572 27620 14600
rect 27614 14560 27620 14572
rect 27672 14560 27678 14612
rect 27798 14600 27804 14612
rect 27759 14572 27804 14600
rect 27798 14560 27804 14572
rect 27856 14560 27862 14612
rect 30006 14600 30012 14612
rect 29967 14572 30012 14600
rect 30006 14560 30012 14572
rect 30064 14560 30070 14612
rect 32582 14600 32588 14612
rect 32543 14572 32588 14600
rect 32582 14560 32588 14572
rect 32640 14560 32646 14612
rect 32950 14560 32956 14612
rect 33008 14600 33014 14612
rect 33045 14603 33103 14609
rect 33045 14600 33057 14603
rect 33008 14572 33057 14600
rect 33008 14560 33014 14572
rect 33045 14569 33057 14572
rect 33091 14569 33103 14603
rect 33045 14563 33103 14569
rect 35253 14603 35311 14609
rect 35253 14569 35265 14603
rect 35299 14600 35311 14603
rect 35526 14600 35532 14612
rect 35299 14572 35532 14600
rect 35299 14569 35311 14572
rect 35253 14563 35311 14569
rect 35526 14560 35532 14572
rect 35584 14560 35590 14612
rect 37274 14600 37280 14612
rect 37235 14572 37280 14600
rect 37274 14560 37280 14572
rect 37332 14560 37338 14612
rect 19426 14464 19432 14476
rect 19387 14436 19432 14464
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 24118 14464 24124 14476
rect 23952 14436 24124 14464
rect 21542 14396 21548 14408
rect 21503 14368 21548 14396
rect 21542 14356 21548 14368
rect 21600 14356 21606 14408
rect 21634 14396 21692 14402
rect 21913 14399 21971 14405
rect 21634 14362 21646 14396
rect 21680 14362 21692 14396
rect 21634 14356 21692 14362
rect 21729 14393 21787 14399
rect 21729 14359 21741 14393
rect 21775 14359 21787 14393
rect 21913 14365 21925 14399
rect 21959 14365 21971 14399
rect 21913 14359 21971 14365
rect 19696 14331 19754 14337
rect 19696 14297 19708 14331
rect 19742 14328 19754 14331
rect 20438 14328 20444 14340
rect 19742 14300 20444 14328
rect 19742 14297 19754 14300
rect 19696 14291 19754 14297
rect 20438 14288 20444 14300
rect 20496 14288 20502 14340
rect 21358 14328 21364 14340
rect 20548 14300 21364 14328
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20548 14260 20576 14300
rect 21358 14288 21364 14300
rect 21416 14328 21422 14340
rect 21649 14328 21677 14356
rect 21729 14353 21787 14359
rect 21416 14300 21677 14328
rect 21416 14288 21422 14300
rect 20806 14260 20812 14272
rect 20128 14232 20576 14260
rect 20767 14232 20812 14260
rect 20128 14220 20134 14232
rect 20806 14220 20812 14232
rect 20864 14220 20870 14272
rect 21266 14220 21272 14272
rect 21324 14260 21330 14272
rect 21744 14260 21772 14353
rect 21324 14232 21772 14260
rect 21928 14260 21956 14359
rect 23566 14356 23572 14408
rect 23624 14362 23630 14408
rect 23661 14399 23719 14405
rect 23850 14399 23908 14405
rect 23661 14365 23673 14399
rect 23707 14365 23719 14399
rect 23661 14362 23719 14365
rect 23624 14359 23719 14362
rect 23750 14393 23808 14399
rect 23750 14359 23762 14393
rect 23796 14362 23808 14393
rect 23850 14365 23862 14399
rect 23896 14396 23908 14399
rect 23952 14396 23980 14436
rect 24118 14424 24124 14436
rect 24176 14424 24182 14476
rect 24670 14424 24676 14476
rect 24728 14464 24734 14476
rect 24949 14467 25007 14473
rect 24949 14464 24961 14467
rect 24728 14436 24961 14464
rect 24728 14424 24734 14436
rect 24949 14433 24961 14436
rect 24995 14433 25007 14467
rect 24949 14427 25007 14433
rect 28718 14424 28724 14476
rect 28776 14464 28782 14476
rect 31205 14467 31263 14473
rect 31205 14464 31217 14467
rect 28776 14436 31217 14464
rect 28776 14424 28782 14436
rect 31205 14433 31217 14436
rect 31251 14433 31263 14467
rect 32600 14464 32628 14560
rect 32600 14436 33272 14464
rect 31205 14427 31263 14433
rect 23896 14368 23980 14396
rect 24029 14399 24087 14405
rect 23896 14365 23908 14368
rect 23796 14359 23809 14362
rect 23850 14359 23908 14365
rect 24029 14365 24041 14399
rect 24075 14396 24087 14399
rect 25774 14396 25780 14408
rect 24075 14368 25780 14396
rect 24075 14365 24087 14368
rect 24029 14359 24087 14365
rect 23624 14356 23704 14359
rect 23584 14334 23704 14356
rect 23750 14353 23809 14359
rect 23768 14334 23809 14353
rect 23781 14328 23809 14334
rect 23934 14328 23940 14340
rect 23781 14300 23940 14328
rect 23934 14288 23940 14300
rect 23992 14288 23998 14340
rect 24044 14260 24072 14359
rect 25774 14356 25780 14368
rect 25832 14356 25838 14408
rect 27982 14356 27988 14408
rect 28040 14396 28046 14408
rect 28445 14399 28503 14405
rect 28445 14396 28457 14399
rect 28040 14368 28457 14396
rect 28040 14356 28046 14368
rect 28445 14365 28457 14368
rect 28491 14365 28503 14399
rect 28445 14359 28503 14365
rect 28629 14399 28687 14405
rect 28629 14365 28641 14399
rect 28675 14365 28687 14399
rect 30190 14396 30196 14408
rect 30151 14368 30196 14396
rect 28629 14359 28687 14365
rect 25222 14337 25228 14340
rect 25216 14291 25228 14337
rect 25280 14328 25286 14340
rect 27433 14331 27491 14337
rect 25280 14300 25316 14328
rect 25222 14288 25228 14291
rect 25280 14288 25286 14300
rect 27433 14297 27445 14331
rect 27479 14328 27491 14331
rect 27522 14328 27528 14340
rect 27479 14300 27528 14328
rect 27479 14297 27491 14300
rect 27433 14291 27491 14297
rect 27522 14288 27528 14300
rect 27580 14288 27586 14340
rect 27706 14337 27712 14340
rect 27649 14331 27712 14337
rect 27649 14297 27661 14331
rect 27695 14297 27712 14331
rect 27649 14291 27712 14297
rect 27706 14288 27712 14291
rect 27764 14288 27770 14340
rect 27890 14288 27896 14340
rect 27948 14328 27954 14340
rect 28644 14328 28672 14359
rect 30190 14356 30196 14368
rect 30248 14356 30254 14408
rect 30650 14356 30656 14408
rect 30708 14396 30714 14408
rect 31461 14399 31519 14405
rect 31461 14396 31473 14399
rect 30708 14368 31473 14396
rect 30708 14356 30714 14368
rect 31461 14365 31473 14368
rect 31507 14365 31519 14399
rect 33042 14396 33048 14408
rect 33003 14368 33048 14396
rect 31461 14359 31519 14365
rect 33042 14356 33048 14368
rect 33100 14356 33106 14408
rect 33244 14405 33272 14436
rect 35894 14424 35900 14476
rect 35952 14464 35958 14476
rect 35952 14436 35997 14464
rect 35952 14424 35958 14436
rect 33229 14399 33287 14405
rect 33229 14365 33241 14399
rect 33275 14365 33287 14399
rect 35434 14396 35440 14408
rect 35395 14368 35440 14396
rect 33229 14359 33287 14365
rect 35434 14356 35440 14368
rect 35492 14356 35498 14408
rect 36164 14399 36222 14405
rect 36164 14365 36176 14399
rect 36210 14396 36222 14399
rect 37458 14396 37464 14408
rect 36210 14368 37464 14396
rect 36210 14365 36222 14368
rect 36164 14359 36222 14365
rect 37458 14356 37464 14368
rect 37516 14356 37522 14408
rect 28902 14328 28908 14340
rect 27948 14300 28908 14328
rect 27948 14288 27954 14300
rect 28902 14288 28908 14300
rect 28960 14288 28966 14340
rect 26326 14260 26332 14272
rect 21928 14232 24072 14260
rect 26287 14232 26332 14260
rect 21324 14220 21330 14232
rect 26326 14220 26332 14232
rect 26384 14220 26390 14272
rect 28629 14263 28687 14269
rect 28629 14229 28641 14263
rect 28675 14260 28687 14263
rect 28994 14260 29000 14272
rect 28675 14232 29000 14260
rect 28675 14229 28687 14232
rect 28629 14223 28687 14229
rect 28994 14220 29000 14232
rect 29052 14220 29058 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 20438 14056 20444 14068
rect 19803 14028 20300 14056
rect 20399 14028 20444 14056
rect 19803 13988 19831 14028
rect 19720 13960 19831 13988
rect 20272 13988 20300 14028
rect 20438 14016 20444 14028
rect 20496 14016 20502 14068
rect 22922 14056 22928 14068
rect 22883 14028 22928 14056
rect 22922 14016 22928 14028
rect 22980 14016 22986 14068
rect 24029 14059 24087 14065
rect 24029 14025 24041 14059
rect 24075 14056 24087 14059
rect 24118 14056 24124 14068
rect 24075 14028 24124 14056
rect 24075 14025 24087 14028
rect 24029 14019 24087 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 25133 14059 25191 14065
rect 25133 14025 25145 14059
rect 25179 14056 25191 14059
rect 25222 14056 25228 14068
rect 25179 14028 25228 14056
rect 25179 14025 25191 14028
rect 25133 14019 25191 14025
rect 25222 14016 25228 14028
rect 25280 14016 25286 14068
rect 27890 14056 27896 14068
rect 25516 14028 27896 14056
rect 20272 13960 21036 13988
rect 18877 13923 18935 13929
rect 18877 13889 18889 13923
rect 18923 13920 18935 13923
rect 19518 13920 19524 13932
rect 18923 13892 19524 13920
rect 18923 13889 18935 13892
rect 18877 13883 18935 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19720 13929 19748 13960
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 19886 13920 19892 13932
rect 19847 13892 19892 13920
rect 19705 13883 19763 13889
rect 19886 13880 19892 13892
rect 19944 13880 19950 13932
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13889 20039 13923
rect 19981 13883 20039 13889
rect 18969 13855 19027 13861
rect 18969 13821 18981 13855
rect 19015 13852 19027 13855
rect 19426 13852 19432 13864
rect 19015 13824 19432 13852
rect 19015 13821 19027 13824
rect 18969 13815 19027 13821
rect 19426 13812 19432 13824
rect 19484 13812 19490 13864
rect 19996 13852 20024 13883
rect 20070 13880 20076 13932
rect 20128 13920 20134 13932
rect 20268 13923 20326 13929
rect 20128 13892 20173 13920
rect 20128 13880 20134 13892
rect 20268 13889 20280 13923
rect 20314 13920 20326 13923
rect 20438 13920 20444 13932
rect 20314 13892 20444 13920
rect 20314 13889 20326 13892
rect 20268 13883 20326 13889
rect 20438 13880 20444 13892
rect 20496 13880 20502 13932
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20772 13892 20913 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 21008 13920 21036 13960
rect 21358 13948 21364 14000
rect 21416 13988 21422 14000
rect 23934 13988 23940 14000
rect 21416 13960 23940 13988
rect 21416 13948 21422 13960
rect 22186 13920 22192 13932
rect 21008 13892 22192 13920
rect 20901 13883 20959 13889
rect 22186 13880 22192 13892
rect 22244 13880 22250 13932
rect 22370 13920 22376 13932
rect 22331 13892 22376 13920
rect 22370 13880 22376 13892
rect 22428 13880 22434 13932
rect 22572 13929 22600 13960
rect 23934 13948 23940 13960
rect 23992 13988 23998 14000
rect 25516 13988 25544 14028
rect 27890 14016 27896 14028
rect 27948 14016 27954 14068
rect 30193 14059 30251 14065
rect 30193 14056 30205 14059
rect 28644 14028 30205 14056
rect 23992 13960 25544 13988
rect 23992 13948 23998 13960
rect 22557 13923 22615 13929
rect 22557 13889 22569 13923
rect 22603 13889 22615 13923
rect 22738 13920 22744 13932
rect 22699 13892 22744 13920
rect 22557 13883 22615 13889
rect 22738 13880 22744 13892
rect 22796 13880 22802 13932
rect 23750 13920 23756 13932
rect 23711 13892 23756 13920
rect 23750 13880 23756 13892
rect 23808 13880 23814 13932
rect 25516 13929 25544 13960
rect 26418 13948 26424 14000
rect 26476 13988 26482 14000
rect 27709 13991 27767 13997
rect 26476 13960 27660 13988
rect 26476 13948 26482 13960
rect 25409 13923 25467 13929
rect 25409 13889 25421 13923
rect 25455 13889 25467 13923
rect 25409 13883 25467 13889
rect 25501 13923 25559 13929
rect 25501 13889 25513 13923
rect 25547 13889 25559 13923
rect 25501 13883 25559 13889
rect 19996 13824 21128 13852
rect 21100 13793 21128 13824
rect 21174 13812 21180 13864
rect 21232 13852 21238 13864
rect 22002 13852 22008 13864
rect 21232 13824 22008 13852
rect 21232 13812 21238 13824
rect 22002 13812 22008 13824
rect 22060 13852 22066 13864
rect 22462 13852 22468 13864
rect 22060 13824 22324 13852
rect 22423 13824 22468 13852
rect 22060 13812 22066 13824
rect 20993 13787 21051 13793
rect 20993 13784 21005 13787
rect 20272 13756 21005 13784
rect 19153 13719 19211 13725
rect 19153 13685 19165 13719
rect 19199 13716 19211 13719
rect 19794 13716 19800 13728
rect 19199 13688 19800 13716
rect 19199 13685 19211 13688
rect 19153 13679 19211 13685
rect 19794 13676 19800 13688
rect 19852 13716 19858 13728
rect 20272 13716 20300 13756
rect 20993 13753 21005 13756
rect 21039 13753 21051 13787
rect 20993 13747 21051 13753
rect 21085 13787 21143 13793
rect 21085 13753 21097 13787
rect 21131 13753 21143 13787
rect 22296 13784 22324 13824
rect 22462 13812 22468 13824
rect 22520 13812 22526 13864
rect 24029 13855 24087 13861
rect 24029 13821 24041 13855
rect 24075 13852 24087 13855
rect 24854 13852 24860 13864
rect 24075 13824 24860 13852
rect 24075 13821 24087 13824
rect 24029 13815 24087 13821
rect 24044 13784 24072 13815
rect 24854 13812 24860 13824
rect 24912 13812 24918 13864
rect 25424 13852 25452 13883
rect 25590 13880 25596 13932
rect 25648 13920 25654 13932
rect 25648 13892 25693 13920
rect 25648 13880 25654 13892
rect 25774 13880 25780 13932
rect 25832 13920 25838 13932
rect 27632 13920 27660 13960
rect 27709 13957 27721 13991
rect 27755 13988 27767 13991
rect 28074 13988 28080 14000
rect 27755 13960 28080 13988
rect 27755 13957 27767 13960
rect 27709 13951 27767 13957
rect 28074 13948 28080 13960
rect 28132 13948 28138 14000
rect 28644 13932 28672 14028
rect 30193 14025 30205 14028
rect 30239 14025 30251 14059
rect 30193 14019 30251 14025
rect 35434 14016 35440 14068
rect 35492 14056 35498 14068
rect 36173 14059 36231 14065
rect 36173 14056 36185 14059
rect 35492 14028 36185 14056
rect 35492 14016 35498 14028
rect 36173 14025 36185 14028
rect 36219 14025 36231 14059
rect 36173 14019 36231 14025
rect 29178 13988 29184 14000
rect 28966 13960 29184 13988
rect 27893 13923 27951 13929
rect 27893 13920 27905 13923
rect 25832 13892 26464 13920
rect 27632 13892 27905 13920
rect 25832 13880 25838 13892
rect 26326 13852 26332 13864
rect 25424 13824 26332 13852
rect 26326 13812 26332 13824
rect 26384 13812 26390 13864
rect 26436 13852 26464 13892
rect 27893 13889 27905 13892
rect 27939 13920 27951 13923
rect 28626 13920 28632 13932
rect 27939 13892 28632 13920
rect 27939 13889 27951 13892
rect 27893 13883 27951 13889
rect 28626 13880 28632 13892
rect 28684 13880 28690 13932
rect 28718 13880 28724 13932
rect 28776 13920 28782 13932
rect 28813 13923 28871 13929
rect 28813 13920 28825 13923
rect 28776 13892 28825 13920
rect 28776 13880 28782 13892
rect 28813 13889 28825 13892
rect 28859 13889 28871 13923
rect 28966 13920 28994 13960
rect 29178 13948 29184 13960
rect 29236 13948 29242 14000
rect 29086 13929 29092 13932
rect 28813 13883 28871 13889
rect 28920 13892 28994 13920
rect 28920 13852 28948 13892
rect 29080 13883 29092 13929
rect 29144 13920 29150 13932
rect 35989 13923 36047 13929
rect 29144 13892 29180 13920
rect 29086 13880 29092 13883
rect 29144 13880 29150 13892
rect 35989 13889 36001 13923
rect 36035 13920 36047 13923
rect 38102 13920 38108 13932
rect 36035 13892 38108 13920
rect 36035 13889 36047 13892
rect 35989 13883 36047 13889
rect 38102 13880 38108 13892
rect 38160 13880 38166 13932
rect 35802 13852 35808 13864
rect 26436 13824 28948 13852
rect 35763 13824 35808 13852
rect 35802 13812 35808 13824
rect 35860 13812 35866 13864
rect 22296 13756 24072 13784
rect 21085 13747 21143 13753
rect 23842 13716 23848 13728
rect 19852 13688 20300 13716
rect 23803 13688 23848 13716
rect 19852 13676 19858 13688
rect 23842 13676 23848 13688
rect 23900 13676 23906 13728
rect 28077 13719 28135 13725
rect 28077 13685 28089 13719
rect 28123 13716 28135 13719
rect 28350 13716 28356 13728
rect 28123 13688 28356 13716
rect 28123 13685 28135 13688
rect 28077 13679 28135 13685
rect 28350 13676 28356 13688
rect 28408 13676 28414 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 19886 13472 19892 13524
rect 19944 13512 19950 13524
rect 19981 13515 20039 13521
rect 19981 13512 19993 13515
rect 19944 13484 19993 13512
rect 19944 13472 19950 13484
rect 19981 13481 19993 13484
rect 20027 13481 20039 13515
rect 19981 13475 20039 13481
rect 20533 13515 20591 13521
rect 20533 13481 20545 13515
rect 20579 13512 20591 13515
rect 20622 13512 20628 13524
rect 20579 13484 20628 13512
rect 20579 13481 20591 13484
rect 20533 13475 20591 13481
rect 19518 13404 19524 13456
rect 19576 13444 19582 13456
rect 20548 13444 20576 13475
rect 20622 13472 20628 13484
rect 20680 13472 20686 13524
rect 21266 13512 21272 13524
rect 21227 13484 21272 13512
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 22462 13472 22468 13524
rect 22520 13512 22526 13524
rect 23017 13515 23075 13521
rect 23017 13512 23029 13515
rect 22520 13484 23029 13512
rect 22520 13472 22526 13484
rect 23017 13481 23029 13484
rect 23063 13481 23075 13515
rect 23017 13475 23075 13481
rect 24949 13515 25007 13521
rect 24949 13481 24961 13515
rect 24995 13512 25007 13515
rect 25590 13512 25596 13524
rect 24995 13484 25596 13512
rect 24995 13481 25007 13484
rect 24949 13475 25007 13481
rect 25590 13472 25596 13484
rect 25648 13472 25654 13524
rect 28537 13515 28595 13521
rect 28537 13481 28549 13515
rect 28583 13512 28595 13515
rect 29086 13512 29092 13524
rect 28583 13484 29092 13512
rect 28583 13481 28595 13484
rect 28537 13475 28595 13481
rect 29086 13472 29092 13484
rect 29144 13472 29150 13524
rect 30101 13515 30159 13521
rect 30101 13481 30113 13515
rect 30147 13512 30159 13515
rect 30190 13512 30196 13524
rect 30147 13484 30196 13512
rect 30147 13481 30159 13484
rect 30101 13475 30159 13481
rect 30190 13472 30196 13484
rect 30248 13472 30254 13524
rect 27338 13444 27344 13456
rect 19576 13416 20576 13444
rect 26712 13416 27344 13444
rect 19576 13404 19582 13416
rect 19613 13379 19671 13385
rect 19613 13345 19625 13379
rect 19659 13376 19671 13379
rect 20714 13376 20720 13388
rect 19659 13348 20720 13376
rect 19659 13345 19671 13348
rect 19613 13339 19671 13345
rect 20714 13336 20720 13348
rect 20772 13336 20778 13388
rect 22094 13336 22100 13388
rect 22152 13376 22158 13388
rect 22373 13379 22431 13385
rect 22373 13376 22385 13379
rect 22152 13348 22385 13376
rect 22152 13336 22158 13348
rect 22373 13345 22385 13348
rect 22419 13345 22431 13379
rect 22373 13339 22431 13345
rect 24673 13379 24731 13385
rect 24673 13345 24685 13379
rect 24719 13376 24731 13379
rect 26237 13379 26295 13385
rect 26237 13376 26249 13379
rect 24719 13348 26249 13376
rect 24719 13345 24731 13348
rect 24673 13339 24731 13345
rect 26237 13345 26249 13348
rect 26283 13345 26295 13379
rect 26237 13339 26295 13345
rect 26712 13320 26740 13416
rect 27338 13404 27344 13416
rect 27396 13444 27402 13456
rect 27982 13444 27988 13456
rect 27396 13416 27660 13444
rect 27943 13416 27988 13444
rect 27396 13404 27402 13416
rect 26973 13379 27031 13385
rect 26973 13345 26985 13379
rect 27019 13376 27031 13379
rect 27430 13376 27436 13388
rect 27019 13348 27436 13376
rect 27019 13345 27031 13348
rect 26973 13339 27031 13345
rect 27430 13336 27436 13348
rect 27488 13336 27494 13388
rect 19794 13308 19800 13320
rect 19755 13280 19800 13308
rect 19794 13268 19800 13280
rect 19852 13268 19858 13320
rect 20438 13308 20444 13320
rect 20351 13280 20444 13308
rect 20438 13268 20444 13280
rect 20496 13308 20502 13320
rect 20806 13308 20812 13320
rect 20496 13280 20812 13308
rect 20496 13268 20502 13280
rect 20806 13268 20812 13280
rect 20864 13268 20870 13320
rect 20898 13268 20904 13320
rect 20956 13308 20962 13320
rect 21177 13311 21235 13317
rect 21177 13308 21189 13311
rect 20956 13280 21189 13308
rect 20956 13268 20962 13280
rect 21177 13277 21189 13280
rect 21223 13277 21235 13311
rect 21358 13308 21364 13320
rect 21319 13280 21364 13308
rect 21177 13271 21235 13277
rect 21358 13268 21364 13280
rect 21416 13268 21422 13320
rect 22462 13268 22468 13320
rect 22520 13308 22526 13320
rect 22741 13311 22799 13317
rect 22741 13308 22753 13311
rect 22520 13280 22753 13308
rect 22520 13268 22526 13280
rect 22741 13277 22753 13280
rect 22787 13277 22799 13311
rect 22741 13271 22799 13277
rect 22833 13311 22891 13317
rect 22833 13277 22845 13311
rect 22879 13308 22891 13311
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 22879 13280 23489 13308
rect 22879 13277 22891 13280
rect 22833 13271 22891 13277
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 23661 13311 23719 13317
rect 23661 13277 23673 13311
rect 23707 13308 23719 13311
rect 23842 13308 23848 13320
rect 23707 13280 23848 13308
rect 23707 13277 23719 13280
rect 23661 13271 23719 13277
rect 22278 13200 22284 13252
rect 22336 13240 22342 13252
rect 22848 13240 22876 13271
rect 22336 13212 22876 13240
rect 23676 13240 23704 13271
rect 23842 13268 23848 13280
rect 23900 13268 23906 13320
rect 23934 13268 23940 13320
rect 23992 13308 23998 13320
rect 24949 13311 25007 13317
rect 23992 13280 24037 13308
rect 23992 13268 23998 13280
rect 24949 13277 24961 13311
rect 24995 13277 25007 13311
rect 24949 13271 25007 13277
rect 25133 13311 25191 13317
rect 25133 13277 25145 13311
rect 25179 13308 25191 13311
rect 25958 13308 25964 13320
rect 25179 13280 25964 13308
rect 25179 13277 25191 13280
rect 25133 13271 25191 13277
rect 24670 13240 24676 13252
rect 23676 13212 24676 13240
rect 22336 13200 22342 13212
rect 24670 13200 24676 13212
rect 24728 13200 24734 13252
rect 24964 13240 24992 13271
rect 25958 13268 25964 13280
rect 26016 13268 26022 13320
rect 26053 13311 26111 13317
rect 26053 13277 26065 13311
rect 26099 13277 26111 13311
rect 26694 13308 26700 13320
rect 26607 13280 26700 13308
rect 26053 13271 26111 13277
rect 26068 13240 26096 13271
rect 26694 13268 26700 13280
rect 26752 13268 26758 13320
rect 26786 13268 26792 13320
rect 26844 13308 26850 13320
rect 27632 13317 27660 13416
rect 27982 13404 27988 13416
rect 28040 13404 28046 13456
rect 28994 13404 29000 13456
rect 29052 13444 29058 13456
rect 29052 13416 29132 13444
rect 29052 13404 29058 13416
rect 27709 13379 27767 13385
rect 27709 13345 27721 13379
rect 27755 13345 27767 13379
rect 27709 13339 27767 13345
rect 27617 13311 27675 13317
rect 26844 13280 27476 13308
rect 26844 13268 26850 13280
rect 26973 13243 27031 13249
rect 26973 13240 26985 13243
rect 24964 13212 26985 13240
rect 26973 13209 26985 13212
rect 27019 13209 27031 13243
rect 27448 13240 27476 13280
rect 27617 13277 27629 13311
rect 27663 13277 27675 13311
rect 27617 13271 27675 13277
rect 27724 13240 27752 13339
rect 28626 13268 28632 13320
rect 28684 13308 28690 13320
rect 28767 13311 28825 13317
rect 28767 13308 28779 13311
rect 28684 13280 28779 13308
rect 28684 13268 28690 13280
rect 28767 13277 28779 13280
rect 28813 13277 28825 13311
rect 28902 13308 28908 13320
rect 28863 13280 28908 13308
rect 28767 13271 28825 13277
rect 28902 13268 28908 13280
rect 28960 13268 28966 13320
rect 29018 13311 29076 13317
rect 29018 13277 29030 13311
rect 29064 13308 29076 13311
rect 29104 13308 29132 13416
rect 29733 13379 29791 13385
rect 29733 13345 29745 13379
rect 29779 13376 29791 13379
rect 32766 13376 32772 13388
rect 29779 13348 32772 13376
rect 29779 13345 29791 13348
rect 29733 13339 29791 13345
rect 32766 13336 32772 13348
rect 32824 13376 32830 13388
rect 35802 13376 35808 13388
rect 32824 13348 35808 13376
rect 32824 13336 32830 13348
rect 35802 13336 35808 13348
rect 35860 13336 35866 13388
rect 29064 13280 29132 13308
rect 29064 13277 29076 13280
rect 29018 13271 29076 13277
rect 29178 13268 29184 13320
rect 29236 13308 29242 13320
rect 29236 13280 29281 13308
rect 29236 13268 29242 13280
rect 29638 13268 29644 13320
rect 29696 13308 29702 13320
rect 29917 13311 29975 13317
rect 29917 13308 29929 13311
rect 29696 13280 29929 13308
rect 29696 13268 29702 13280
rect 29917 13277 29929 13280
rect 29963 13277 29975 13311
rect 29917 13271 29975 13277
rect 28258 13240 28264 13252
rect 27448 13212 28264 13240
rect 26973 13203 27031 13209
rect 28258 13200 28264 13212
rect 28316 13200 28322 13252
rect 23658 13132 23664 13184
rect 23716 13172 23722 13184
rect 23845 13175 23903 13181
rect 23845 13172 23857 13175
rect 23716 13144 23857 13172
rect 23716 13132 23722 13144
rect 23845 13141 23857 13144
rect 23891 13141 23903 13175
rect 23845 13135 23903 13141
rect 24854 13132 24860 13184
rect 24912 13172 24918 13184
rect 25593 13175 25651 13181
rect 25593 13172 25605 13175
rect 24912 13144 25605 13172
rect 24912 13132 24918 13144
rect 25593 13141 25605 13144
rect 25639 13172 25651 13175
rect 27246 13172 27252 13184
rect 25639 13144 27252 13172
rect 25639 13141 25651 13144
rect 25593 13135 25651 13141
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 20073 12971 20131 12977
rect 20073 12937 20085 12971
rect 20119 12968 20131 12971
rect 20714 12968 20720 12980
rect 20119 12940 20720 12968
rect 20119 12937 20131 12940
rect 20073 12931 20131 12937
rect 20714 12928 20720 12940
rect 20772 12928 20778 12980
rect 22370 12968 22376 12980
rect 22331 12940 22376 12968
rect 22370 12928 22376 12940
rect 22428 12928 22434 12980
rect 23750 12928 23756 12980
rect 23808 12968 23814 12980
rect 24121 12971 24179 12977
rect 24121 12968 24133 12971
rect 23808 12940 24133 12968
rect 23808 12928 23814 12940
rect 24121 12937 24133 12940
rect 24167 12937 24179 12971
rect 24670 12968 24676 12980
rect 24631 12940 24676 12968
rect 24121 12931 24179 12937
rect 24670 12928 24676 12940
rect 24728 12928 24734 12980
rect 28258 12968 28264 12980
rect 28219 12940 28264 12968
rect 28258 12928 28264 12940
rect 28316 12928 28322 12980
rect 27341 12903 27399 12909
rect 27341 12869 27353 12903
rect 27387 12900 27399 12903
rect 28074 12900 28080 12912
rect 27387 12872 28080 12900
rect 27387 12869 27399 12872
rect 27341 12863 27399 12869
rect 28074 12860 28080 12872
rect 28132 12860 28138 12912
rect 20254 12832 20260 12844
rect 20215 12804 20260 12832
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 22278 12832 22284 12844
rect 22239 12804 22284 12832
rect 22278 12792 22284 12804
rect 22336 12792 22342 12844
rect 22462 12832 22468 12844
rect 22423 12804 22468 12832
rect 22462 12792 22468 12804
rect 22520 12792 22526 12844
rect 22738 12792 22744 12844
rect 22796 12832 22802 12844
rect 22925 12835 22983 12841
rect 22925 12832 22937 12835
rect 22796 12804 22937 12832
rect 22796 12792 22802 12804
rect 22925 12801 22937 12804
rect 22971 12801 22983 12835
rect 22925 12795 22983 12801
rect 23017 12835 23075 12841
rect 23017 12801 23029 12835
rect 23063 12832 23075 12835
rect 23658 12832 23664 12844
rect 23063 12804 23664 12832
rect 23063 12801 23075 12804
rect 23017 12795 23075 12801
rect 23658 12792 23664 12804
rect 23716 12792 23722 12844
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12832 23995 12835
rect 24026 12832 24032 12844
rect 23983 12804 24032 12832
rect 23983 12801 23995 12804
rect 23937 12795 23995 12801
rect 24026 12792 24032 12804
rect 24084 12832 24090 12844
rect 24581 12835 24639 12841
rect 24581 12832 24593 12835
rect 24084 12804 24593 12832
rect 24084 12792 24090 12804
rect 24581 12801 24593 12804
rect 24627 12801 24639 12835
rect 24762 12832 24768 12844
rect 24581 12795 24639 12801
rect 24688 12804 24768 12832
rect 20530 12764 20536 12776
rect 20491 12736 20536 12764
rect 20530 12724 20536 12736
rect 20588 12724 20594 12776
rect 23201 12767 23259 12773
rect 23201 12733 23213 12767
rect 23247 12764 23259 12767
rect 23247 12736 23281 12764
rect 23247 12733 23259 12736
rect 23201 12727 23259 12733
rect 22094 12656 22100 12708
rect 22152 12696 22158 12708
rect 23216 12696 23244 12727
rect 23382 12724 23388 12776
rect 23440 12764 23446 12776
rect 23753 12767 23811 12773
rect 23753 12764 23765 12767
rect 23440 12736 23765 12764
rect 23440 12724 23446 12736
rect 23753 12733 23765 12736
rect 23799 12764 23811 12767
rect 24688 12764 24716 12804
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 25409 12835 25467 12841
rect 25409 12801 25421 12835
rect 25455 12832 25467 12835
rect 26237 12835 26295 12841
rect 26237 12832 26249 12835
rect 25455 12804 26249 12832
rect 25455 12801 25467 12804
rect 25409 12795 25467 12801
rect 26237 12801 26249 12804
rect 26283 12832 26295 12835
rect 26326 12832 26332 12844
rect 26283 12804 26332 12832
rect 26283 12801 26295 12804
rect 26237 12795 26295 12801
rect 26326 12792 26332 12804
rect 26384 12792 26390 12844
rect 27430 12792 27436 12844
rect 27488 12832 27494 12844
rect 28169 12835 28227 12841
rect 28169 12832 28181 12835
rect 27488 12804 28181 12832
rect 27488 12792 27494 12804
rect 28169 12801 28181 12804
rect 28215 12801 28227 12835
rect 28350 12832 28356 12844
rect 28311 12804 28356 12832
rect 28169 12795 28227 12801
rect 28350 12792 28356 12804
rect 28408 12792 28414 12844
rect 23799 12736 24716 12764
rect 25317 12767 25375 12773
rect 23799 12733 23811 12736
rect 23753 12727 23811 12733
rect 25317 12733 25329 12767
rect 25363 12764 25375 12767
rect 26513 12767 26571 12773
rect 26513 12764 26525 12767
rect 25363 12736 26525 12764
rect 25363 12733 25375 12736
rect 25317 12727 25375 12733
rect 26513 12733 26525 12736
rect 26559 12764 26571 12767
rect 27246 12764 27252 12776
rect 26559 12736 27252 12764
rect 26559 12733 26571 12736
rect 26513 12727 26571 12733
rect 23934 12696 23940 12708
rect 22152 12668 23940 12696
rect 22152 12656 22158 12668
rect 23934 12656 23940 12668
rect 23992 12696 23998 12708
rect 25332 12696 25360 12727
rect 27246 12724 27252 12736
rect 27304 12764 27310 12776
rect 27617 12767 27675 12773
rect 27617 12764 27629 12767
rect 27304 12736 27629 12764
rect 27304 12724 27310 12736
rect 27617 12733 27629 12736
rect 27663 12733 27675 12767
rect 27617 12727 27675 12733
rect 23992 12668 25360 12696
rect 25777 12699 25835 12705
rect 23992 12656 23998 12668
rect 25777 12665 25789 12699
rect 25823 12696 25835 12699
rect 26234 12696 26240 12708
rect 25823 12668 26240 12696
rect 25823 12665 25835 12668
rect 25777 12659 25835 12665
rect 26234 12656 26240 12668
rect 26292 12656 26298 12708
rect 26326 12656 26332 12708
rect 26384 12696 26390 12708
rect 26384 12668 26429 12696
rect 26384 12656 26390 12668
rect 20438 12628 20444 12640
rect 20399 12600 20444 12628
rect 20438 12588 20444 12600
rect 20496 12588 20502 12640
rect 23109 12631 23167 12637
rect 23109 12597 23121 12631
rect 23155 12628 23167 12631
rect 23474 12628 23480 12640
rect 23155 12600 23480 12628
rect 23155 12597 23167 12600
rect 23109 12591 23167 12597
rect 23474 12588 23480 12600
rect 23532 12588 23538 12640
rect 26418 12588 26424 12640
rect 26476 12628 26482 12640
rect 26476 12600 26521 12628
rect 26476 12588 26482 12600
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 19797 12427 19855 12433
rect 19797 12393 19809 12427
rect 19843 12424 19855 12427
rect 20254 12424 20260 12436
rect 19843 12396 20260 12424
rect 19843 12393 19855 12396
rect 19797 12387 19855 12393
rect 20254 12384 20260 12396
rect 20312 12384 20318 12436
rect 20530 12384 20536 12436
rect 20588 12424 20594 12436
rect 21361 12427 21419 12433
rect 21361 12424 21373 12427
rect 20588 12396 21373 12424
rect 20588 12384 20594 12396
rect 21361 12393 21373 12396
rect 21407 12393 21419 12427
rect 23017 12427 23075 12433
rect 23017 12424 23029 12427
rect 21361 12387 21419 12393
rect 21468 12396 23029 12424
rect 20898 12356 20904 12368
rect 20859 12328 20904 12356
rect 20898 12316 20904 12328
rect 20956 12316 20962 12368
rect 21468 12356 21496 12396
rect 23017 12393 23029 12396
rect 23063 12393 23075 12427
rect 23017 12387 23075 12393
rect 24762 12384 24768 12436
rect 24820 12424 24826 12436
rect 25961 12427 26019 12433
rect 25961 12424 25973 12427
rect 24820 12396 25973 12424
rect 24820 12384 24826 12396
rect 25961 12393 25973 12396
rect 26007 12393 26019 12427
rect 27338 12424 27344 12436
rect 27299 12396 27344 12424
rect 25961 12387 26019 12393
rect 27338 12384 27344 12396
rect 27396 12384 27402 12436
rect 21284 12328 21496 12356
rect 19720 12260 20392 12288
rect 19426 12180 19432 12232
rect 19484 12220 19490 12232
rect 19720 12229 19748 12260
rect 19705 12223 19763 12229
rect 19705 12220 19717 12223
rect 19484 12192 19717 12220
rect 19484 12180 19490 12192
rect 19705 12189 19717 12192
rect 19751 12189 19763 12223
rect 19705 12183 19763 12189
rect 19889 12223 19947 12229
rect 19889 12189 19901 12223
rect 19935 12189 19947 12223
rect 19889 12183 19947 12189
rect 19904 12084 19932 12183
rect 20364 12152 20392 12260
rect 20438 12248 20444 12300
rect 20496 12288 20502 12300
rect 20625 12291 20683 12297
rect 20625 12288 20637 12291
rect 20496 12260 20637 12288
rect 20496 12248 20502 12260
rect 20625 12257 20637 12260
rect 20671 12288 20683 12291
rect 21284 12288 21312 12328
rect 22462 12316 22468 12368
rect 22520 12356 22526 12368
rect 22557 12359 22615 12365
rect 22557 12356 22569 12359
rect 22520 12328 22569 12356
rect 22520 12316 22526 12328
rect 22557 12325 22569 12328
rect 22603 12325 22615 12359
rect 22557 12319 22615 12325
rect 23293 12359 23351 12365
rect 23293 12325 23305 12359
rect 23339 12356 23351 12359
rect 24026 12356 24032 12368
rect 23339 12328 24032 12356
rect 23339 12325 23351 12328
rect 23293 12319 23351 12325
rect 22094 12288 22100 12300
rect 20671 12260 21312 12288
rect 21376 12260 22100 12288
rect 20671 12257 20683 12260
rect 20625 12251 20683 12257
rect 20533 12223 20591 12229
rect 20533 12189 20545 12223
rect 20579 12220 20591 12223
rect 20806 12220 20812 12232
rect 20579 12192 20812 12220
rect 20579 12189 20591 12192
rect 20533 12183 20591 12189
rect 20806 12180 20812 12192
rect 20864 12180 20870 12232
rect 21376 12229 21404 12260
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 22572 12288 22600 12319
rect 24026 12316 24032 12328
rect 24084 12316 24090 12368
rect 26234 12316 26240 12368
rect 26292 12356 26298 12368
rect 26329 12359 26387 12365
rect 26329 12356 26341 12359
rect 26292 12328 26341 12356
rect 26292 12316 26298 12328
rect 26329 12325 26341 12328
rect 26375 12325 26387 12359
rect 26329 12319 26387 12325
rect 26510 12316 26516 12368
rect 26568 12356 26574 12368
rect 26568 12328 27476 12356
rect 26568 12316 26574 12328
rect 23385 12291 23443 12297
rect 23385 12288 23397 12291
rect 22572 12260 23397 12288
rect 23385 12257 23397 12260
rect 23431 12257 23443 12291
rect 26786 12288 26792 12300
rect 23385 12251 23443 12257
rect 26252 12260 26792 12288
rect 21361 12223 21419 12229
rect 21361 12220 21373 12223
rect 21192 12192 21373 12220
rect 21192 12152 21220 12192
rect 21361 12189 21373 12192
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21545 12223 21603 12229
rect 21545 12220 21557 12223
rect 21508 12192 21557 12220
rect 21508 12180 21514 12192
rect 21545 12189 21557 12192
rect 21591 12189 21603 12223
rect 21545 12183 21603 12189
rect 22189 12223 22247 12229
rect 22189 12189 22201 12223
rect 22235 12220 22247 12223
rect 22738 12220 22744 12232
rect 22235 12192 22744 12220
rect 22235 12189 22247 12192
rect 22189 12183 22247 12189
rect 22738 12180 22744 12192
rect 22796 12180 22802 12232
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12220 23259 12223
rect 23290 12220 23296 12232
rect 23247 12192 23296 12220
rect 23247 12189 23259 12192
rect 23201 12183 23259 12189
rect 23290 12180 23296 12192
rect 23348 12180 23354 12232
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 26252 12229 26280 12260
rect 26786 12248 26792 12260
rect 26844 12248 26850 12300
rect 26145 12223 26203 12229
rect 23532 12192 23577 12220
rect 23532 12180 23538 12192
rect 26145 12189 26157 12223
rect 26191 12189 26203 12223
rect 26145 12183 26203 12189
rect 26237 12223 26295 12229
rect 26237 12189 26249 12223
rect 26283 12189 26295 12223
rect 26237 12183 26295 12189
rect 20364 12124 21220 12152
rect 21468 12084 21496 12180
rect 26160 12152 26188 12183
rect 26418 12180 26424 12232
rect 26476 12220 26482 12232
rect 27246 12220 27252 12232
rect 26476 12192 26521 12220
rect 27207 12192 27252 12220
rect 26476 12180 26482 12192
rect 27246 12180 27252 12192
rect 27304 12180 27310 12232
rect 27448 12229 27476 12328
rect 27433 12223 27491 12229
rect 27433 12189 27445 12223
rect 27479 12189 27491 12223
rect 27433 12183 27491 12189
rect 26694 12152 26700 12164
rect 26160 12124 26700 12152
rect 26694 12112 26700 12124
rect 26752 12112 26758 12164
rect 19904 12056 21496 12084
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 20806 11880 20812 11892
rect 20767 11852 20812 11880
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 24026 11880 24032 11892
rect 23987 11852 24032 11880
rect 24026 11840 24032 11852
rect 24084 11840 24090 11892
rect 20254 11704 20260 11756
rect 20312 11744 20318 11756
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 20312 11716 20361 11744
rect 20312 11704 20318 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 23658 11744 23664 11756
rect 23619 11716 23664 11744
rect 20349 11707 20407 11713
rect 23658 11704 23664 11716
rect 23716 11704 23722 11756
rect 23753 11679 23811 11685
rect 23753 11645 23765 11679
rect 23799 11676 23811 11679
rect 23934 11676 23940 11688
rect 23799 11648 23940 11676
rect 23799 11645 23811 11648
rect 23753 11639 23811 11645
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 20530 11540 20536 11552
rect 20491 11512 20536 11540
rect 20530 11500 20536 11512
rect 20588 11500 20594 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1762 10452 1768 10464
rect 1723 10424 1768 10452
rect 1762 10412 1768 10424
rect 1820 10412 1826 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 29914 8916 29920 8968
rect 29972 8956 29978 8968
rect 38013 8959 38071 8965
rect 38013 8956 38025 8959
rect 29972 8928 38025 8956
rect 29972 8916 29978 8928
rect 38013 8925 38025 8928
rect 38059 8925 38071 8959
rect 38013 8919 38071 8925
rect 38194 8820 38200 8832
rect 38155 8792 38200 8820
rect 38194 8780 38200 8792
rect 38252 8780 38258 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 29638 2592 29644 2644
rect 29696 2632 29702 2644
rect 29733 2635 29791 2641
rect 29733 2632 29745 2635
rect 29696 2604 29745 2632
rect 29696 2592 29702 2604
rect 29733 2601 29745 2604
rect 29779 2601 29791 2635
rect 38102 2632 38108 2644
rect 38063 2604 38108 2632
rect 29733 2595 29791 2601
rect 38102 2592 38108 2604
rect 38160 2592 38166 2644
rect 1854 2496 1860 2508
rect 1815 2468 1860 2496
rect 1854 2456 1860 2468
rect 1912 2456 1918 2508
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1581 2431 1639 2437
rect 1581 2428 1593 2431
rect 72 2400 1593 2428
rect 72 2388 78 2400
rect 1581 2397 1593 2400
rect 1627 2397 1639 2431
rect 1581 2391 1639 2397
rect 9674 2388 9680 2440
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 9953 2391 10011 2397
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 28994 2388 29000 2440
rect 29052 2428 29058 2440
rect 29917 2431 29975 2437
rect 29917 2428 29929 2431
rect 29052 2400 29929 2428
rect 29052 2388 29058 2400
rect 29917 2397 29929 2400
rect 29963 2397 29975 2431
rect 29917 2391 29975 2397
rect 38289 2431 38347 2437
rect 38289 2397 38301 2431
rect 38335 2428 38347 2431
rect 38654 2428 38660 2440
rect 38335 2400 38660 2428
rect 38335 2397 38347 2400
rect 38289 2391 38347 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19613 2295 19671 2301
rect 19613 2292 19625 2295
rect 19392 2264 19625 2292
rect 19392 2252 19398 2264
rect 19613 2261 19625 2264
rect 19659 2261 19671 2295
rect 19613 2255 19671 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 29644 37408 29696 37460
rect 39304 37408 39356 37460
rect 664 37204 716 37256
rect 10324 37204 10376 37256
rect 19984 37204 20036 37256
rect 32312 37204 32364 37256
rect 1584 37111 1636 37120
rect 1584 37077 1593 37111
rect 1593 37077 1627 37111
rect 1627 37077 1636 37111
rect 1584 37068 1636 37077
rect 10600 37111 10652 37120
rect 10600 37077 10609 37111
rect 10609 37077 10643 37111
rect 10643 37077 10652 37111
rect 10600 37068 10652 37077
rect 24492 37068 24544 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 32312 36907 32364 36916
rect 32312 36873 32321 36907
rect 32321 36873 32355 36907
rect 32355 36873 32364 36907
rect 32312 36864 32364 36873
rect 32496 36771 32548 36780
rect 32496 36737 32505 36771
rect 32505 36737 32539 36771
rect 32539 36737 32548 36771
rect 32496 36728 32548 36737
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 26976 34076 27028 34128
rect 31208 34076 31260 34128
rect 26792 34051 26844 34060
rect 26792 34017 26801 34051
rect 26801 34017 26835 34051
rect 26835 34017 26844 34051
rect 26792 34008 26844 34017
rect 25136 33940 25188 33992
rect 26516 33983 26568 33992
rect 26516 33949 26525 33983
rect 26525 33949 26559 33983
rect 26559 33949 26568 33983
rect 26516 33940 26568 33949
rect 27620 33983 27672 33992
rect 27620 33949 27629 33983
rect 27629 33949 27663 33983
rect 27663 33949 27672 33983
rect 27620 33940 27672 33949
rect 24860 33872 24912 33924
rect 28264 33940 28316 33992
rect 28540 33983 28592 33992
rect 28540 33949 28549 33983
rect 28549 33949 28583 33983
rect 28583 33949 28592 33983
rect 28540 33940 28592 33949
rect 29184 33983 29236 33992
rect 29184 33949 29193 33983
rect 29193 33949 29227 33983
rect 29227 33949 29236 33983
rect 29184 33940 29236 33949
rect 30104 33940 30156 33992
rect 31024 33983 31076 33992
rect 30196 33872 30248 33924
rect 31024 33949 31033 33983
rect 31033 33949 31067 33983
rect 31067 33949 31076 33983
rect 31024 33940 31076 33949
rect 31668 33940 31720 33992
rect 23848 33804 23900 33856
rect 28356 33804 28408 33856
rect 28448 33804 28500 33856
rect 30564 33804 30616 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 26516 33643 26568 33652
rect 26516 33609 26525 33643
rect 26525 33609 26559 33643
rect 26559 33609 26568 33643
rect 26516 33600 26568 33609
rect 27620 33600 27672 33652
rect 30104 33600 30156 33652
rect 24032 33464 24084 33516
rect 24860 33507 24912 33516
rect 24860 33473 24869 33507
rect 24869 33473 24903 33507
rect 24903 33473 24912 33507
rect 24860 33464 24912 33473
rect 27252 33464 27304 33516
rect 27620 33507 27672 33516
rect 27620 33473 27629 33507
rect 27629 33473 27663 33507
rect 27663 33473 27672 33507
rect 27620 33464 27672 33473
rect 30380 33532 30432 33584
rect 30104 33507 30156 33516
rect 23940 33439 23992 33448
rect 23940 33405 23949 33439
rect 23949 33405 23983 33439
rect 23983 33405 23992 33439
rect 23940 33396 23992 33405
rect 26056 33439 26108 33448
rect 26056 33405 26065 33439
rect 26065 33405 26099 33439
rect 26099 33405 26108 33439
rect 26056 33396 26108 33405
rect 28448 33439 28500 33448
rect 28448 33405 28457 33439
rect 28457 33405 28491 33439
rect 28491 33405 28500 33439
rect 28448 33396 28500 33405
rect 30104 33473 30113 33507
rect 30113 33473 30147 33507
rect 30147 33473 30156 33507
rect 30104 33464 30156 33473
rect 30196 33464 30248 33516
rect 30564 33507 30616 33516
rect 30564 33473 30573 33507
rect 30573 33473 30607 33507
rect 30607 33473 30616 33507
rect 30564 33464 30616 33473
rect 34520 33396 34572 33448
rect 23480 33328 23532 33380
rect 25136 33328 25188 33380
rect 26516 33260 26568 33312
rect 29092 33328 29144 33380
rect 34152 33328 34204 33380
rect 28908 33260 28960 33312
rect 30564 33260 30616 33312
rect 31392 33303 31444 33312
rect 31392 33269 31401 33303
rect 31401 33269 31435 33303
rect 31435 33269 31444 33303
rect 31392 33260 31444 33269
rect 33968 33303 34020 33312
rect 33968 33269 33977 33303
rect 33977 33269 34011 33303
rect 34011 33269 34020 33303
rect 33968 33260 34020 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 26792 33056 26844 33108
rect 27620 33056 27672 33108
rect 29184 33099 29236 33108
rect 29184 33065 29193 33099
rect 29193 33065 29227 33099
rect 29227 33065 29236 33099
rect 29184 33056 29236 33065
rect 30564 33056 30616 33108
rect 31392 33056 31444 33108
rect 33968 33099 34020 33108
rect 33968 33065 33977 33099
rect 33977 33065 34011 33099
rect 34011 33065 34020 33099
rect 33968 33056 34020 33065
rect 23480 32988 23532 33040
rect 23756 33031 23808 33040
rect 23756 32997 23765 33031
rect 23765 32997 23799 33031
rect 23799 32997 23808 33031
rect 23756 32988 23808 32997
rect 24860 32988 24912 33040
rect 24584 32920 24636 32972
rect 34520 32988 34572 33040
rect 28264 32920 28316 32972
rect 28908 32920 28960 32972
rect 29736 32920 29788 32972
rect 34060 32963 34112 32972
rect 34060 32929 34069 32963
rect 34069 32929 34103 32963
rect 34103 32929 34112 32963
rect 34060 32920 34112 32929
rect 23848 32852 23900 32904
rect 23940 32852 23992 32904
rect 24860 32852 24912 32904
rect 25136 32895 25188 32904
rect 25136 32861 25145 32895
rect 25145 32861 25179 32895
rect 25179 32861 25188 32895
rect 25136 32852 25188 32861
rect 25228 32852 25280 32904
rect 25964 32852 26016 32904
rect 26976 32895 27028 32904
rect 26976 32861 26985 32895
rect 26985 32861 27019 32895
rect 27019 32861 27028 32895
rect 26976 32852 27028 32861
rect 27252 32852 27304 32904
rect 31208 32895 31260 32904
rect 25044 32784 25096 32836
rect 31208 32861 31217 32895
rect 31217 32861 31251 32895
rect 31251 32861 31260 32895
rect 31208 32852 31260 32861
rect 33692 32895 33744 32904
rect 33692 32861 33701 32895
rect 33701 32861 33735 32895
rect 33735 32861 33744 32895
rect 33692 32852 33744 32861
rect 33784 32895 33836 32904
rect 33784 32861 33793 32895
rect 33793 32861 33827 32895
rect 33827 32861 33836 32895
rect 33784 32852 33836 32861
rect 28448 32784 28500 32836
rect 30380 32827 30432 32836
rect 30380 32793 30389 32827
rect 30389 32793 30423 32827
rect 30423 32793 30432 32827
rect 30380 32784 30432 32793
rect 30564 32827 30616 32836
rect 30564 32793 30573 32827
rect 30573 32793 30607 32827
rect 30607 32793 30616 32827
rect 30564 32784 30616 32793
rect 34152 32784 34204 32836
rect 24032 32716 24084 32768
rect 24952 32759 25004 32768
rect 24952 32725 24961 32759
rect 24961 32725 24995 32759
rect 24995 32725 25004 32759
rect 24952 32716 25004 32725
rect 26516 32716 26568 32768
rect 30840 32716 30892 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 25228 32555 25280 32564
rect 25228 32521 25237 32555
rect 25237 32521 25271 32555
rect 25271 32521 25280 32555
rect 25228 32512 25280 32521
rect 25964 32555 26016 32564
rect 25964 32521 25973 32555
rect 25973 32521 26007 32555
rect 26007 32521 26016 32555
rect 25964 32512 26016 32521
rect 25136 32376 25188 32428
rect 25780 32376 25832 32428
rect 28172 32376 28224 32428
rect 28448 32512 28500 32564
rect 30380 32512 30432 32564
rect 31024 32512 31076 32564
rect 28632 32419 28684 32428
rect 23756 32351 23808 32360
rect 23756 32317 23765 32351
rect 23765 32317 23799 32351
rect 23799 32317 23808 32351
rect 23756 32308 23808 32317
rect 24216 32283 24268 32292
rect 24216 32249 24225 32283
rect 24225 32249 24259 32283
rect 24259 32249 24268 32283
rect 24216 32240 24268 32249
rect 24860 32240 24912 32292
rect 26148 32308 26200 32360
rect 27620 32308 27672 32360
rect 28632 32385 28641 32419
rect 28641 32385 28675 32419
rect 28675 32385 28684 32419
rect 28632 32376 28684 32385
rect 29092 32419 29144 32428
rect 29092 32385 29101 32419
rect 29101 32385 29135 32419
rect 29135 32385 29144 32419
rect 29092 32376 29144 32385
rect 30564 32419 30616 32428
rect 25228 32240 25280 32292
rect 21272 32172 21324 32224
rect 24400 32172 24452 32224
rect 24768 32172 24820 32224
rect 25780 32215 25832 32224
rect 25780 32181 25789 32215
rect 25789 32181 25823 32215
rect 25823 32181 25832 32215
rect 25780 32172 25832 32181
rect 28080 32172 28132 32224
rect 28540 32240 28592 32292
rect 30564 32385 30573 32419
rect 30573 32385 30607 32419
rect 30607 32385 30616 32419
rect 30564 32376 30616 32385
rect 30840 32376 30892 32428
rect 30932 32419 30984 32428
rect 30932 32385 30941 32419
rect 30941 32385 30975 32419
rect 30975 32385 30984 32419
rect 33784 32512 33836 32564
rect 30932 32376 30984 32385
rect 33876 32376 33928 32428
rect 34060 32376 34112 32428
rect 37648 32419 37700 32428
rect 31668 32308 31720 32360
rect 34428 32351 34480 32360
rect 34428 32317 34437 32351
rect 34437 32317 34471 32351
rect 34471 32317 34480 32351
rect 34428 32308 34480 32317
rect 37648 32385 37657 32419
rect 37657 32385 37691 32419
rect 37691 32385 37700 32419
rect 37648 32376 37700 32385
rect 36268 32308 36320 32360
rect 28632 32172 28684 32224
rect 30932 32240 30984 32292
rect 33692 32240 33744 32292
rect 30748 32172 30800 32224
rect 37188 32172 37240 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 31668 31968 31720 32020
rect 31760 31968 31812 32020
rect 34428 31968 34480 32020
rect 36268 32011 36320 32020
rect 36268 31977 36277 32011
rect 36277 31977 36311 32011
rect 36311 31977 36320 32011
rect 36268 31968 36320 31977
rect 24032 31900 24084 31952
rect 24768 31900 24820 31952
rect 21272 31875 21324 31884
rect 21272 31841 21281 31875
rect 21281 31841 21315 31875
rect 21315 31841 21324 31875
rect 21272 31832 21324 31841
rect 21364 31832 21416 31884
rect 1584 31764 1636 31816
rect 27252 31900 27304 31952
rect 27436 31943 27488 31952
rect 27436 31909 27445 31943
rect 27445 31909 27479 31943
rect 27479 31909 27488 31943
rect 27436 31900 27488 31909
rect 25044 31807 25096 31816
rect 25044 31773 25053 31807
rect 25053 31773 25087 31807
rect 25087 31773 25096 31807
rect 25228 31807 25280 31816
rect 25044 31764 25096 31773
rect 25228 31773 25237 31807
rect 25237 31773 25271 31807
rect 25271 31773 25280 31807
rect 25228 31764 25280 31773
rect 26056 31807 26108 31816
rect 26056 31773 26065 31807
rect 26065 31773 26099 31807
rect 26099 31773 26108 31807
rect 26056 31764 26108 31773
rect 37280 31900 37332 31952
rect 26608 31696 26660 31748
rect 26240 31628 26292 31680
rect 27620 31696 27672 31748
rect 28356 31807 28408 31816
rect 28356 31773 28365 31807
rect 28365 31773 28399 31807
rect 28399 31773 28408 31807
rect 28356 31764 28408 31773
rect 28632 31764 28684 31816
rect 29736 31807 29788 31816
rect 29736 31773 29745 31807
rect 29745 31773 29779 31807
rect 29779 31773 29788 31807
rect 29736 31764 29788 31773
rect 28908 31628 28960 31680
rect 30288 31696 30340 31748
rect 30748 31764 30800 31816
rect 32496 31807 32548 31816
rect 32496 31773 32505 31807
rect 32505 31773 32539 31807
rect 32539 31773 32548 31807
rect 32496 31764 32548 31773
rect 34612 31764 34664 31816
rect 32404 31696 32456 31748
rect 35532 31764 35584 31816
rect 36912 31807 36964 31816
rect 36912 31773 36921 31807
rect 36921 31773 36955 31807
rect 36955 31773 36964 31807
rect 36912 31764 36964 31773
rect 37832 31764 37884 31816
rect 38292 31807 38344 31816
rect 38292 31773 38301 31807
rect 38301 31773 38335 31807
rect 38335 31773 38344 31807
rect 38292 31764 38344 31773
rect 30104 31628 30156 31680
rect 36728 31671 36780 31680
rect 36728 31637 36737 31671
rect 36737 31637 36771 31671
rect 36771 31637 36780 31671
rect 36728 31628 36780 31637
rect 37464 31671 37516 31680
rect 37464 31637 37473 31671
rect 37473 31637 37507 31671
rect 37507 31637 37516 31671
rect 37464 31628 37516 31637
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 26240 31424 26292 31476
rect 27620 31424 27672 31476
rect 30196 31424 30248 31476
rect 32404 31467 32456 31476
rect 32404 31433 32413 31467
rect 32413 31433 32447 31467
rect 32447 31433 32456 31467
rect 32404 31424 32456 31433
rect 37648 31424 37700 31476
rect 28080 31399 28132 31408
rect 28080 31365 28114 31399
rect 28114 31365 28132 31399
rect 28080 31356 28132 31365
rect 20076 31288 20128 31340
rect 22928 31288 22980 31340
rect 26056 31288 26108 31340
rect 27160 31288 27212 31340
rect 30288 31356 30340 31408
rect 29736 31288 29788 31340
rect 31668 31331 31720 31340
rect 31668 31297 31677 31331
rect 31677 31297 31711 31331
rect 31711 31297 31720 31331
rect 31668 31288 31720 31297
rect 36728 31356 36780 31408
rect 33232 31331 33284 31340
rect 33232 31297 33241 31331
rect 33241 31297 33275 31331
rect 33275 31297 33284 31331
rect 33232 31288 33284 31297
rect 35532 31331 35584 31340
rect 35532 31297 35541 31331
rect 35541 31297 35575 31331
rect 35575 31297 35584 31331
rect 35532 31288 35584 31297
rect 36176 31288 36228 31340
rect 19432 31220 19484 31272
rect 22836 31220 22888 31272
rect 34428 31220 34480 31272
rect 20260 31084 20312 31136
rect 21732 31084 21784 31136
rect 22376 31127 22428 31136
rect 22376 31093 22385 31127
rect 22385 31093 22419 31127
rect 22419 31093 22428 31127
rect 22376 31084 22428 31093
rect 28448 31084 28500 31136
rect 31300 31084 31352 31136
rect 37372 31084 37424 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 17408 30880 17460 30932
rect 20352 30880 20404 30932
rect 22468 30880 22520 30932
rect 22836 30923 22888 30932
rect 22836 30889 22845 30923
rect 22845 30889 22879 30923
rect 22879 30889 22888 30923
rect 22836 30880 22888 30889
rect 24952 30880 25004 30932
rect 25504 30880 25556 30932
rect 29736 30923 29788 30932
rect 29736 30889 29745 30923
rect 29745 30889 29779 30923
rect 29779 30889 29788 30923
rect 29736 30880 29788 30889
rect 30104 30923 30156 30932
rect 30104 30889 30113 30923
rect 30113 30889 30147 30923
rect 30147 30889 30156 30923
rect 30104 30880 30156 30889
rect 33232 30880 33284 30932
rect 36176 30880 36228 30932
rect 36912 30880 36964 30932
rect 29368 30812 29420 30864
rect 35532 30812 35584 30864
rect 25780 30787 25832 30796
rect 25780 30753 25789 30787
rect 25789 30753 25823 30787
rect 25823 30753 25832 30787
rect 25780 30744 25832 30753
rect 36912 30787 36964 30796
rect 1584 30719 1636 30728
rect 1584 30685 1593 30719
rect 1593 30685 1627 30719
rect 1627 30685 1636 30719
rect 1584 30676 1636 30685
rect 17040 30719 17092 30728
rect 17040 30685 17049 30719
rect 17049 30685 17083 30719
rect 17083 30685 17092 30719
rect 17040 30676 17092 30685
rect 18604 30676 18656 30728
rect 20260 30719 20312 30728
rect 20260 30685 20269 30719
rect 20269 30685 20303 30719
rect 20303 30685 20312 30719
rect 20260 30676 20312 30685
rect 21364 30676 21416 30728
rect 22008 30676 22060 30728
rect 24584 30719 24636 30728
rect 24584 30685 24593 30719
rect 24593 30685 24627 30719
rect 24627 30685 24636 30719
rect 24584 30676 24636 30685
rect 25044 30676 25096 30728
rect 26240 30719 26292 30728
rect 20168 30608 20220 30660
rect 21732 30651 21784 30660
rect 21732 30617 21766 30651
rect 21766 30617 21784 30651
rect 21732 30608 21784 30617
rect 26240 30685 26249 30719
rect 26249 30685 26283 30719
rect 26283 30685 26292 30719
rect 26240 30676 26292 30685
rect 26608 30676 26660 30728
rect 26884 30719 26936 30728
rect 26884 30685 26893 30719
rect 26893 30685 26927 30719
rect 26927 30685 26936 30719
rect 26884 30676 26936 30685
rect 27620 30676 27672 30728
rect 29184 30719 29236 30728
rect 29184 30685 29193 30719
rect 29193 30685 29227 30719
rect 29227 30685 29236 30719
rect 29184 30676 29236 30685
rect 29644 30676 29696 30728
rect 36912 30753 36921 30787
rect 36921 30753 36955 30787
rect 36955 30753 36964 30787
rect 36912 30744 36964 30753
rect 30196 30719 30248 30728
rect 30196 30685 30205 30719
rect 30205 30685 30239 30719
rect 30239 30685 30248 30719
rect 30196 30676 30248 30685
rect 30288 30676 30340 30728
rect 25872 30608 25924 30660
rect 28724 30608 28776 30660
rect 29000 30608 29052 30660
rect 32496 30676 32548 30728
rect 35716 30676 35768 30728
rect 36176 30719 36228 30728
rect 31300 30651 31352 30660
rect 1768 30583 1820 30592
rect 1768 30549 1777 30583
rect 1777 30549 1811 30583
rect 1811 30549 1820 30583
rect 1768 30540 1820 30549
rect 17224 30540 17276 30592
rect 19340 30540 19392 30592
rect 20352 30583 20404 30592
rect 20352 30549 20361 30583
rect 20361 30549 20395 30583
rect 20395 30549 20404 30583
rect 20352 30540 20404 30549
rect 24860 30540 24912 30592
rect 27252 30540 27304 30592
rect 28816 30540 28868 30592
rect 31300 30617 31334 30651
rect 31334 30617 31352 30651
rect 31300 30608 31352 30617
rect 31392 30608 31444 30660
rect 33968 30608 34020 30660
rect 36176 30685 36185 30719
rect 36185 30685 36219 30719
rect 36219 30685 36228 30719
rect 36176 30676 36228 30685
rect 37188 30719 37240 30728
rect 37188 30685 37222 30719
rect 37222 30685 37240 30719
rect 37188 30676 37240 30685
rect 36268 30608 36320 30660
rect 31852 30540 31904 30592
rect 34060 30540 34112 30592
rect 35624 30540 35676 30592
rect 37924 30540 37976 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 19616 30336 19668 30388
rect 20260 30336 20312 30388
rect 17132 30243 17184 30252
rect 16580 30132 16632 30184
rect 17132 30209 17141 30243
rect 17141 30209 17175 30243
rect 17175 30209 17184 30243
rect 17132 30200 17184 30209
rect 18512 30200 18564 30252
rect 19340 30268 19392 30320
rect 19524 30268 19576 30320
rect 22008 30268 22060 30320
rect 28724 30336 28776 30388
rect 29184 30336 29236 30388
rect 33968 30379 34020 30388
rect 33968 30345 33977 30379
rect 33977 30345 34011 30379
rect 34011 30345 34020 30379
rect 33968 30336 34020 30345
rect 35532 30336 35584 30388
rect 18880 30175 18932 30184
rect 18880 30141 18889 30175
rect 18889 30141 18923 30175
rect 18923 30141 18932 30175
rect 18880 30132 18932 30141
rect 19064 30132 19116 30184
rect 19432 30200 19484 30252
rect 19892 30200 19944 30252
rect 22468 30243 22520 30252
rect 22468 30209 22477 30243
rect 22477 30209 22511 30243
rect 22511 30209 22520 30243
rect 22468 30200 22520 30209
rect 22836 30243 22888 30252
rect 22836 30209 22845 30243
rect 22845 30209 22879 30243
rect 22879 30209 22888 30243
rect 22836 30200 22888 30209
rect 19616 30132 19668 30184
rect 21916 30132 21968 30184
rect 22192 30175 22244 30184
rect 22192 30141 22201 30175
rect 22201 30141 22235 30175
rect 22235 30141 22244 30175
rect 22192 30132 22244 30141
rect 23480 30132 23532 30184
rect 26240 30268 26292 30320
rect 24952 30200 25004 30252
rect 26056 30200 26108 30252
rect 28908 30268 28960 30320
rect 33692 30268 33744 30320
rect 26608 30243 26660 30252
rect 26608 30209 26617 30243
rect 26617 30209 26651 30243
rect 26651 30209 26660 30243
rect 26608 30200 26660 30209
rect 26976 30200 27028 30252
rect 27160 30243 27212 30252
rect 27160 30209 27169 30243
rect 27169 30209 27203 30243
rect 27203 30209 27212 30243
rect 27160 30200 27212 30209
rect 27436 30243 27488 30252
rect 27436 30209 27470 30243
rect 27470 30209 27488 30243
rect 29368 30243 29420 30252
rect 27436 30200 27488 30209
rect 29368 30209 29377 30243
rect 29377 30209 29411 30243
rect 29411 30209 29420 30243
rect 29368 30200 29420 30209
rect 34152 30243 34204 30252
rect 34152 30209 34161 30243
rect 34161 30209 34195 30243
rect 34195 30209 34204 30243
rect 34152 30200 34204 30209
rect 25504 30175 25556 30184
rect 25504 30141 25513 30175
rect 25513 30141 25547 30175
rect 25547 30141 25556 30175
rect 25504 30132 25556 30141
rect 25780 30132 25832 30184
rect 29460 30175 29512 30184
rect 29460 30141 29469 30175
rect 29469 30141 29503 30175
rect 29503 30141 29512 30175
rect 29460 30132 29512 30141
rect 19800 30064 19852 30116
rect 20812 30064 20864 30116
rect 26884 30064 26936 30116
rect 17408 29996 17460 30048
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 20076 29996 20128 30048
rect 21088 29996 21140 30048
rect 25044 29996 25096 30048
rect 26976 29996 27028 30048
rect 30012 30064 30064 30116
rect 28724 29996 28776 30048
rect 34796 30200 34848 30252
rect 35624 30311 35676 30320
rect 35624 30277 35658 30311
rect 35658 30277 35676 30311
rect 35624 30268 35676 30277
rect 36268 30268 36320 30320
rect 37924 30336 37976 30388
rect 37556 30200 37608 30252
rect 34612 30175 34664 30184
rect 34612 30141 34621 30175
rect 34621 30141 34655 30175
rect 34655 30141 34664 30175
rect 34612 30132 34664 30141
rect 37372 30064 37424 30116
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 17040 29792 17092 29844
rect 18880 29792 18932 29844
rect 19524 29792 19576 29844
rect 19800 29792 19852 29844
rect 20352 29792 20404 29844
rect 22192 29792 22244 29844
rect 22928 29835 22980 29844
rect 22928 29801 22937 29835
rect 22937 29801 22971 29835
rect 22971 29801 22980 29835
rect 22928 29792 22980 29801
rect 24860 29835 24912 29844
rect 24860 29801 24869 29835
rect 24869 29801 24903 29835
rect 24903 29801 24912 29835
rect 24860 29792 24912 29801
rect 24952 29835 25004 29844
rect 24952 29801 24961 29835
rect 24961 29801 24995 29835
rect 24995 29801 25004 29835
rect 25872 29835 25924 29844
rect 24952 29792 25004 29801
rect 25872 29801 25881 29835
rect 25881 29801 25915 29835
rect 25915 29801 25924 29835
rect 25872 29792 25924 29801
rect 26056 29835 26108 29844
rect 26056 29801 26065 29835
rect 26065 29801 26099 29835
rect 26099 29801 26108 29835
rect 26056 29792 26108 29801
rect 27436 29792 27488 29844
rect 29460 29792 29512 29844
rect 34152 29792 34204 29844
rect 34796 29792 34848 29844
rect 36268 29835 36320 29844
rect 36268 29801 36277 29835
rect 36277 29801 36311 29835
rect 36311 29801 36320 29835
rect 36268 29792 36320 29801
rect 16488 29588 16540 29640
rect 17132 29656 17184 29708
rect 17316 29699 17368 29708
rect 17316 29665 17325 29699
rect 17325 29665 17359 29699
rect 17359 29665 17368 29699
rect 17316 29656 17368 29665
rect 18052 29724 18104 29776
rect 20168 29724 20220 29776
rect 21456 29724 21508 29776
rect 21916 29724 21968 29776
rect 18788 29656 18840 29708
rect 17224 29631 17276 29640
rect 17224 29597 17233 29631
rect 17233 29597 17267 29631
rect 17267 29597 17276 29631
rect 17224 29588 17276 29597
rect 18604 29631 18656 29640
rect 18604 29597 18613 29631
rect 18613 29597 18647 29631
rect 18647 29597 18656 29631
rect 18604 29588 18656 29597
rect 18696 29588 18748 29640
rect 1584 29520 1636 29572
rect 18696 29452 18748 29504
rect 20812 29656 20864 29708
rect 21824 29656 21876 29708
rect 24952 29699 25004 29708
rect 24952 29665 24961 29699
rect 24961 29665 24995 29699
rect 24995 29665 25004 29699
rect 24952 29656 25004 29665
rect 19064 29588 19116 29640
rect 20076 29631 20128 29640
rect 19340 29520 19392 29572
rect 20076 29597 20085 29631
rect 20085 29597 20119 29631
rect 20119 29597 20128 29631
rect 20076 29588 20128 29597
rect 21088 29631 21140 29640
rect 20168 29520 20220 29572
rect 21088 29597 21097 29631
rect 21097 29597 21131 29631
rect 21131 29597 21140 29631
rect 21088 29588 21140 29597
rect 22468 29588 22520 29640
rect 22836 29588 22888 29640
rect 23204 29631 23256 29640
rect 23204 29597 23213 29631
rect 23213 29597 23247 29631
rect 23247 29597 23256 29631
rect 23204 29588 23256 29597
rect 24216 29588 24268 29640
rect 25780 29588 25832 29640
rect 26976 29631 27028 29640
rect 26976 29597 26985 29631
rect 26985 29597 27019 29631
rect 27019 29597 27028 29631
rect 26976 29588 27028 29597
rect 22100 29520 22152 29572
rect 23480 29520 23532 29572
rect 27252 29588 27304 29640
rect 28632 29724 28684 29776
rect 30564 29724 30616 29776
rect 37556 29792 37608 29844
rect 28724 29699 28776 29708
rect 28724 29665 28733 29699
rect 28733 29665 28767 29699
rect 28767 29665 28776 29699
rect 28724 29656 28776 29665
rect 28908 29656 28960 29708
rect 36912 29699 36964 29708
rect 36912 29665 36921 29699
rect 36921 29665 36955 29699
rect 36955 29665 36964 29699
rect 36912 29656 36964 29665
rect 28448 29631 28500 29640
rect 28448 29597 28457 29631
rect 28457 29597 28491 29631
rect 28491 29597 28500 29631
rect 28448 29588 28500 29597
rect 28632 29631 28684 29640
rect 28632 29597 28641 29631
rect 28641 29597 28675 29631
rect 28675 29597 28684 29631
rect 28632 29588 28684 29597
rect 27620 29520 27672 29572
rect 30932 29588 30984 29640
rect 31852 29631 31904 29640
rect 31852 29597 31861 29631
rect 31861 29597 31895 29631
rect 31895 29597 31904 29631
rect 31852 29588 31904 29597
rect 32220 29588 32272 29640
rect 33968 29631 34020 29640
rect 33968 29597 33977 29631
rect 33977 29597 34011 29631
rect 34011 29597 34020 29631
rect 33968 29588 34020 29597
rect 34520 29588 34572 29640
rect 32772 29520 32824 29572
rect 34244 29520 34296 29572
rect 22284 29452 22336 29504
rect 22376 29452 22428 29504
rect 23204 29452 23256 29504
rect 28448 29452 28500 29504
rect 28908 29452 28960 29504
rect 29644 29452 29696 29504
rect 31760 29452 31812 29504
rect 34152 29495 34204 29504
rect 34152 29461 34161 29495
rect 34161 29461 34195 29495
rect 34195 29461 34204 29495
rect 35992 29563 36044 29572
rect 35992 29529 36001 29563
rect 36001 29529 36035 29563
rect 36035 29529 36044 29563
rect 35992 29520 36044 29529
rect 37464 29588 37516 29640
rect 37372 29520 37424 29572
rect 34152 29452 34204 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 18604 29248 18656 29300
rect 20168 29248 20220 29300
rect 18512 29180 18564 29232
rect 19248 29180 19300 29232
rect 20076 29180 20128 29232
rect 17040 29112 17092 29164
rect 17408 29155 17460 29164
rect 17408 29121 17417 29155
rect 17417 29121 17451 29155
rect 17451 29121 17460 29155
rect 17408 29112 17460 29121
rect 18696 29155 18748 29164
rect 18696 29121 18705 29155
rect 18705 29121 18739 29155
rect 18739 29121 18748 29155
rect 18696 29112 18748 29121
rect 19340 29112 19392 29164
rect 23756 29248 23808 29300
rect 25044 29248 25096 29300
rect 27620 29248 27672 29300
rect 28632 29248 28684 29300
rect 30932 29291 30984 29300
rect 30932 29257 30941 29291
rect 30941 29257 30975 29291
rect 30975 29257 30984 29291
rect 30932 29248 30984 29257
rect 34244 29291 34296 29300
rect 34244 29257 34253 29291
rect 34253 29257 34287 29291
rect 34287 29257 34296 29291
rect 34244 29248 34296 29257
rect 35716 29248 35768 29300
rect 37832 29291 37884 29300
rect 37832 29257 37841 29291
rect 37841 29257 37875 29291
rect 37875 29257 37884 29291
rect 37832 29248 37884 29257
rect 22376 29155 22428 29164
rect 22376 29121 22385 29155
rect 22385 29121 22419 29155
rect 22419 29121 22428 29155
rect 22376 29112 22428 29121
rect 25780 29112 25832 29164
rect 26424 29155 26476 29164
rect 19984 29044 20036 29096
rect 22008 29044 22060 29096
rect 26424 29121 26433 29155
rect 26433 29121 26467 29155
rect 26467 29121 26476 29155
rect 26424 29112 26476 29121
rect 28540 29180 28592 29232
rect 27068 29044 27120 29096
rect 28264 29112 28316 29164
rect 29460 29180 29512 29232
rect 29368 29112 29420 29164
rect 30288 29180 30340 29232
rect 34152 29180 34204 29232
rect 34336 29180 34388 29232
rect 29644 29112 29696 29164
rect 31760 29155 31812 29164
rect 31760 29121 31769 29155
rect 31769 29121 31803 29155
rect 31803 29121 31812 29155
rect 31760 29112 31812 29121
rect 32772 29155 32824 29164
rect 32772 29121 32781 29155
rect 32781 29121 32815 29155
rect 32815 29121 32824 29155
rect 32772 29112 32824 29121
rect 32864 29155 32916 29164
rect 32864 29121 32873 29155
rect 32873 29121 32907 29155
rect 32907 29121 32916 29155
rect 32864 29112 32916 29121
rect 33232 29112 33284 29164
rect 28448 29044 28500 29096
rect 28540 29044 28592 29096
rect 35348 29155 35400 29164
rect 35348 29121 35357 29155
rect 35357 29121 35391 29155
rect 35391 29121 35400 29155
rect 35348 29112 35400 29121
rect 35992 29180 36044 29232
rect 34520 29044 34572 29096
rect 37280 29112 37332 29164
rect 37924 29180 37976 29232
rect 37648 29155 37700 29164
rect 37648 29121 37657 29155
rect 37657 29121 37691 29155
rect 37691 29121 37700 29155
rect 37648 29112 37700 29121
rect 17316 29019 17368 29028
rect 17316 28985 17325 29019
rect 17325 28985 17359 29019
rect 17359 28985 17368 29019
rect 17316 28976 17368 28985
rect 27436 28976 27488 29028
rect 33416 28976 33468 29028
rect 33508 28976 33560 29028
rect 23572 28908 23624 28960
rect 25688 28951 25740 28960
rect 25688 28917 25697 28951
rect 25697 28917 25731 28951
rect 25731 28917 25740 28951
rect 25688 28908 25740 28917
rect 27804 28951 27856 28960
rect 27804 28917 27813 28951
rect 27813 28917 27847 28951
rect 27847 28917 27856 28951
rect 27804 28908 27856 28917
rect 31668 28908 31720 28960
rect 33968 28951 34020 28960
rect 33968 28917 33977 28951
rect 33977 28917 34011 28951
rect 34011 28917 34020 28951
rect 33968 28908 34020 28917
rect 36176 28908 36228 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 22284 28747 22336 28756
rect 22284 28713 22293 28747
rect 22293 28713 22327 28747
rect 22327 28713 22336 28747
rect 22284 28704 22336 28713
rect 22652 28704 22704 28756
rect 23204 28704 23256 28756
rect 23756 28747 23808 28756
rect 23756 28713 23765 28747
rect 23765 28713 23799 28747
rect 23799 28713 23808 28747
rect 23756 28704 23808 28713
rect 24400 28704 24452 28756
rect 26424 28747 26476 28756
rect 19892 28500 19944 28552
rect 22744 28636 22796 28688
rect 26424 28713 26433 28747
rect 26433 28713 26467 28747
rect 26467 28713 26476 28747
rect 26424 28704 26476 28713
rect 29276 28636 29328 28688
rect 32312 28704 32364 28756
rect 32772 28747 32824 28756
rect 32772 28713 32781 28747
rect 32781 28713 32815 28747
rect 32815 28713 32824 28747
rect 32772 28704 32824 28713
rect 35532 28704 35584 28756
rect 21916 28568 21968 28620
rect 21824 28543 21876 28552
rect 21824 28509 21831 28543
rect 21831 28509 21876 28543
rect 21824 28500 21876 28509
rect 22192 28500 22244 28552
rect 20168 28432 20220 28484
rect 22652 28432 22704 28484
rect 23112 28500 23164 28552
rect 24860 28568 24912 28620
rect 23572 28543 23624 28552
rect 23572 28509 23581 28543
rect 23581 28509 23615 28543
rect 23615 28509 23624 28543
rect 23572 28500 23624 28509
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 26240 28500 26292 28552
rect 27160 28500 27212 28552
rect 27252 28543 27304 28552
rect 27252 28509 27261 28543
rect 27261 28509 27295 28543
rect 27295 28509 27304 28543
rect 27252 28500 27304 28509
rect 28080 28500 28132 28552
rect 30748 28568 30800 28620
rect 34152 28568 34204 28620
rect 28264 28500 28316 28552
rect 25688 28432 25740 28484
rect 27804 28432 27856 28484
rect 27896 28432 27948 28484
rect 28816 28500 28868 28552
rect 31024 28500 31076 28552
rect 31392 28543 31444 28552
rect 31392 28509 31401 28543
rect 31401 28509 31435 28543
rect 31435 28509 31444 28543
rect 31392 28500 31444 28509
rect 31668 28543 31720 28552
rect 31668 28509 31702 28543
rect 31702 28509 31720 28543
rect 31668 28500 31720 28509
rect 33416 28543 33468 28552
rect 33416 28509 33425 28543
rect 33425 28509 33459 28543
rect 33459 28509 33468 28543
rect 33416 28500 33468 28509
rect 31300 28432 31352 28484
rect 32036 28432 32088 28484
rect 32220 28432 32272 28484
rect 34336 28500 34388 28552
rect 36820 28500 36872 28552
rect 34796 28432 34848 28484
rect 35992 28432 36044 28484
rect 21180 28407 21232 28416
rect 21180 28373 21189 28407
rect 21189 28373 21223 28407
rect 21223 28373 21232 28407
rect 21180 28364 21232 28373
rect 21824 28364 21876 28416
rect 22100 28364 22152 28416
rect 27528 28364 27580 28416
rect 27988 28407 28040 28416
rect 27988 28373 27997 28407
rect 27997 28373 28031 28407
rect 28031 28373 28040 28407
rect 27988 28364 28040 28373
rect 30380 28364 30432 28416
rect 30656 28364 30708 28416
rect 33232 28407 33284 28416
rect 33232 28373 33241 28407
rect 33241 28373 33275 28407
rect 33275 28373 33284 28407
rect 33232 28364 33284 28373
rect 34980 28364 35032 28416
rect 35348 28364 35400 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 10600 28160 10652 28212
rect 20168 28135 20220 28144
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 17132 28024 17184 28033
rect 16580 27820 16632 27872
rect 17684 28024 17736 28076
rect 20168 28101 20177 28135
rect 20177 28101 20211 28135
rect 20211 28101 20220 28135
rect 20168 28092 20220 28101
rect 18420 27999 18472 28008
rect 18420 27965 18429 27999
rect 18429 27965 18463 27999
rect 18463 27965 18472 27999
rect 18420 27956 18472 27965
rect 17592 27820 17644 27872
rect 19340 27820 19392 27872
rect 20628 28067 20680 28076
rect 20628 28033 20637 28067
rect 20637 28033 20671 28067
rect 20671 28033 20680 28067
rect 23112 28092 23164 28144
rect 23664 28160 23716 28212
rect 25780 28203 25832 28212
rect 25780 28169 25789 28203
rect 25789 28169 25823 28203
rect 25823 28169 25832 28203
rect 25780 28160 25832 28169
rect 26424 28160 26476 28212
rect 27068 28160 27120 28212
rect 20628 28024 20680 28033
rect 21180 28024 21232 28076
rect 25044 28092 25096 28144
rect 21456 27956 21508 28008
rect 22652 27956 22704 28008
rect 24492 28024 24544 28076
rect 25964 28067 26016 28076
rect 25964 28033 25973 28067
rect 25973 28033 26007 28067
rect 26007 28033 26016 28067
rect 25964 28024 26016 28033
rect 26332 28024 26384 28076
rect 23572 27956 23624 28008
rect 24124 27956 24176 28008
rect 24400 27999 24452 28008
rect 24400 27965 24409 27999
rect 24409 27965 24443 27999
rect 24443 27965 24452 27999
rect 24400 27956 24452 27965
rect 28080 28160 28132 28212
rect 30656 28160 30708 28212
rect 30748 28160 30800 28212
rect 34152 28160 34204 28212
rect 34796 28203 34848 28212
rect 34796 28169 34805 28203
rect 34805 28169 34839 28203
rect 34839 28169 34848 28203
rect 34796 28160 34848 28169
rect 35992 28203 36044 28212
rect 35992 28169 36001 28203
rect 36001 28169 36035 28203
rect 36035 28169 36044 28203
rect 35992 28160 36044 28169
rect 27896 28092 27948 28144
rect 28356 28135 28408 28144
rect 27988 28067 28040 28076
rect 27988 28033 27997 28067
rect 27997 28033 28031 28067
rect 28031 28033 28040 28067
rect 27988 28024 28040 28033
rect 28356 28101 28365 28135
rect 28365 28101 28399 28135
rect 28399 28101 28408 28135
rect 28356 28092 28408 28101
rect 30932 28092 30984 28144
rect 33232 28092 33284 28144
rect 28264 28067 28316 28076
rect 28264 28033 28273 28067
rect 28273 28033 28307 28067
rect 28307 28033 28316 28067
rect 28264 28024 28316 28033
rect 28448 28067 28500 28076
rect 28448 28033 28462 28067
rect 28462 28033 28496 28067
rect 28496 28033 28500 28067
rect 28448 28024 28500 28033
rect 30012 28067 30064 28076
rect 30012 28033 30022 28067
rect 30022 28033 30056 28067
rect 30056 28033 30064 28067
rect 30012 28024 30064 28033
rect 30196 28067 30248 28076
rect 30196 28033 30205 28067
rect 30205 28033 30239 28067
rect 30239 28033 30248 28067
rect 30196 28024 30248 28033
rect 30380 28067 30432 28076
rect 30380 28033 30394 28067
rect 30394 28033 30428 28067
rect 30428 28033 30432 28067
rect 31024 28067 31076 28076
rect 30380 28024 30432 28033
rect 31024 28033 31033 28067
rect 31033 28033 31067 28067
rect 31067 28033 31076 28067
rect 31024 28024 31076 28033
rect 34336 28067 34388 28076
rect 34336 28033 34345 28067
rect 34345 28033 34379 28067
rect 34379 28033 34388 28067
rect 34336 28024 34388 28033
rect 34980 28067 35032 28076
rect 34980 28033 34989 28067
rect 34989 28033 35023 28067
rect 35023 28033 35032 28067
rect 34980 28024 35032 28033
rect 36176 28067 36228 28076
rect 36176 28033 36185 28067
rect 36185 28033 36219 28067
rect 36219 28033 36228 28067
rect 36176 28024 36228 28033
rect 37556 28024 37608 28076
rect 37648 28067 37700 28076
rect 37648 28033 37657 28067
rect 37657 28033 37691 28067
rect 37691 28033 37700 28067
rect 37648 28024 37700 28033
rect 30472 27956 30524 28008
rect 32036 27956 32088 28008
rect 38016 27956 38068 28008
rect 22100 27888 22152 27940
rect 22560 27888 22612 27940
rect 29184 27888 29236 27940
rect 29276 27888 29328 27940
rect 32220 27888 32272 27940
rect 34612 27888 34664 27940
rect 22284 27863 22336 27872
rect 22284 27829 22293 27863
rect 22293 27829 22327 27863
rect 22327 27829 22336 27863
rect 22284 27820 22336 27829
rect 23112 27820 23164 27872
rect 25964 27820 26016 27872
rect 29552 27820 29604 27872
rect 30932 27820 30984 27872
rect 36728 27820 36780 27872
rect 37464 27820 37516 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 18420 27616 18472 27668
rect 22652 27616 22704 27668
rect 27252 27616 27304 27668
rect 34336 27659 34388 27668
rect 34336 27625 34345 27659
rect 34345 27625 34379 27659
rect 34379 27625 34388 27659
rect 34336 27616 34388 27625
rect 35532 27616 35584 27668
rect 17316 27591 17368 27600
rect 16580 27523 16632 27532
rect 16580 27489 16589 27523
rect 16589 27489 16623 27523
rect 16623 27489 16632 27523
rect 16580 27480 16632 27489
rect 17316 27557 17325 27591
rect 17325 27557 17359 27591
rect 17359 27557 17368 27591
rect 17316 27548 17368 27557
rect 17684 27591 17736 27600
rect 17684 27557 17693 27591
rect 17693 27557 17727 27591
rect 17727 27557 17736 27591
rect 17684 27548 17736 27557
rect 18788 27548 18840 27600
rect 20628 27548 20680 27600
rect 23572 27591 23624 27600
rect 23572 27557 23581 27591
rect 23581 27557 23615 27591
rect 23615 27557 23624 27591
rect 23572 27548 23624 27557
rect 25688 27591 25740 27600
rect 25688 27557 25697 27591
rect 25697 27557 25731 27591
rect 25731 27557 25740 27591
rect 25688 27548 25740 27557
rect 17960 27480 18012 27532
rect 23480 27480 23532 27532
rect 17684 27412 17736 27464
rect 17776 27455 17828 27464
rect 17776 27421 17785 27455
rect 17785 27421 17819 27455
rect 17819 27421 17828 27455
rect 17776 27412 17828 27421
rect 17592 27344 17644 27396
rect 19984 27412 20036 27464
rect 22284 27412 22336 27464
rect 23664 27412 23716 27464
rect 18328 27387 18380 27396
rect 18328 27353 18337 27387
rect 18337 27353 18371 27387
rect 18371 27353 18380 27387
rect 18328 27344 18380 27353
rect 24952 27412 25004 27464
rect 26332 27412 26384 27464
rect 28540 27548 28592 27600
rect 30012 27548 30064 27600
rect 30472 27591 30524 27600
rect 27344 27480 27396 27532
rect 29644 27480 29696 27532
rect 30196 27480 30248 27532
rect 27528 27455 27580 27464
rect 25228 27344 25280 27396
rect 26148 27344 26200 27396
rect 27528 27421 27537 27455
rect 27537 27421 27571 27455
rect 27571 27421 27580 27455
rect 27528 27412 27580 27421
rect 27712 27455 27764 27464
rect 27712 27421 27721 27455
rect 27721 27421 27755 27455
rect 27755 27421 27764 27455
rect 27712 27412 27764 27421
rect 27896 27455 27948 27464
rect 27896 27421 27905 27455
rect 27905 27421 27939 27455
rect 27939 27421 27948 27455
rect 27896 27412 27948 27421
rect 28172 27412 28224 27464
rect 29184 27455 29236 27464
rect 29184 27421 29193 27455
rect 29193 27421 29227 27455
rect 29227 27421 29236 27455
rect 29184 27412 29236 27421
rect 29736 27455 29788 27464
rect 29736 27421 29745 27455
rect 29745 27421 29779 27455
rect 29779 27421 29788 27455
rect 29736 27412 29788 27421
rect 29920 27455 29972 27464
rect 29920 27421 29929 27455
rect 29929 27421 29963 27455
rect 29963 27421 29972 27455
rect 29920 27412 29972 27421
rect 30012 27455 30064 27464
rect 30012 27421 30021 27455
rect 30021 27421 30055 27455
rect 30055 27421 30064 27455
rect 30472 27557 30481 27591
rect 30481 27557 30515 27591
rect 30515 27557 30524 27591
rect 30472 27548 30524 27557
rect 33324 27548 33376 27600
rect 33692 27548 33744 27600
rect 33600 27480 33652 27532
rect 36820 27616 36872 27668
rect 30012 27412 30064 27421
rect 32036 27412 32088 27464
rect 34060 27455 34112 27464
rect 34060 27421 34069 27455
rect 34069 27421 34103 27455
rect 34103 27421 34112 27455
rect 34060 27412 34112 27421
rect 35072 27455 35124 27464
rect 35072 27421 35081 27455
rect 35081 27421 35115 27455
rect 35115 27421 35124 27455
rect 35072 27412 35124 27421
rect 35624 27455 35676 27464
rect 35624 27421 35633 27455
rect 35633 27421 35667 27455
rect 35667 27421 35676 27455
rect 35624 27412 35676 27421
rect 35808 27455 35860 27464
rect 35808 27421 35817 27455
rect 35817 27421 35851 27455
rect 35851 27421 35860 27455
rect 35808 27412 35860 27421
rect 36728 27412 36780 27464
rect 18512 27319 18564 27328
rect 18512 27285 18521 27319
rect 18521 27285 18555 27319
rect 18555 27285 18564 27319
rect 18512 27276 18564 27285
rect 24676 27319 24728 27328
rect 24676 27285 24685 27319
rect 24685 27285 24719 27319
rect 24719 27285 24728 27319
rect 24676 27276 24728 27285
rect 26424 27276 26476 27328
rect 27436 27276 27488 27328
rect 28172 27276 28224 27328
rect 29092 27276 29144 27328
rect 29460 27276 29512 27328
rect 30196 27276 30248 27328
rect 31300 27276 31352 27328
rect 32588 27319 32640 27328
rect 32588 27285 32597 27319
rect 32597 27285 32631 27319
rect 32631 27285 32640 27319
rect 32588 27276 32640 27285
rect 34060 27276 34112 27328
rect 35348 27276 35400 27328
rect 36452 27276 36504 27328
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 17776 27072 17828 27124
rect 22744 27115 22796 27124
rect 22744 27081 22753 27115
rect 22753 27081 22787 27115
rect 22787 27081 22796 27115
rect 22744 27072 22796 27081
rect 26332 27115 26384 27124
rect 26332 27081 26357 27115
rect 26357 27081 26384 27115
rect 26332 27072 26384 27081
rect 27436 27072 27488 27124
rect 29736 27072 29788 27124
rect 30288 27072 30340 27124
rect 30380 27072 30432 27124
rect 31024 27072 31076 27124
rect 32220 27072 32272 27124
rect 32772 27072 32824 27124
rect 35072 27072 35124 27124
rect 35808 27072 35860 27124
rect 24676 27004 24728 27056
rect 26148 27047 26200 27056
rect 26148 27013 26157 27047
rect 26157 27013 26191 27047
rect 26191 27013 26200 27047
rect 26148 27004 26200 27013
rect 27896 27004 27948 27056
rect 17132 26936 17184 26988
rect 17960 26979 18012 26988
rect 17960 26945 17969 26979
rect 17969 26945 18003 26979
rect 18003 26945 18012 26979
rect 17960 26936 18012 26945
rect 18512 26936 18564 26988
rect 17500 26868 17552 26920
rect 17776 26911 17828 26920
rect 17776 26877 17785 26911
rect 17785 26877 17819 26911
rect 17819 26877 17828 26911
rect 17776 26868 17828 26877
rect 19064 26979 19116 26988
rect 19064 26945 19073 26979
rect 19073 26945 19107 26979
rect 19107 26945 19116 26979
rect 19064 26936 19116 26945
rect 19248 26979 19300 26988
rect 19248 26945 19257 26979
rect 19257 26945 19291 26979
rect 19291 26945 19300 26979
rect 19248 26936 19300 26945
rect 18512 26732 18564 26784
rect 19340 26800 19392 26852
rect 22192 26979 22244 26988
rect 22192 26945 22201 26979
rect 22201 26945 22235 26979
rect 22235 26945 22244 26979
rect 22192 26936 22244 26945
rect 22560 26979 22612 26988
rect 22560 26945 22569 26979
rect 22569 26945 22603 26979
rect 22603 26945 22612 26979
rect 22560 26936 22612 26945
rect 28172 26979 28224 26988
rect 28172 26945 28181 26979
rect 28181 26945 28215 26979
rect 28215 26945 28224 26979
rect 28172 26936 28224 26945
rect 28264 26979 28316 26988
rect 28264 26945 28274 26979
rect 28274 26945 28308 26979
rect 28308 26945 28316 26979
rect 28264 26936 28316 26945
rect 22100 26868 22152 26920
rect 21364 26800 21416 26852
rect 22652 26868 22704 26920
rect 19984 26732 20036 26784
rect 21088 26775 21140 26784
rect 21088 26741 21097 26775
rect 21097 26741 21131 26775
rect 21131 26741 21140 26775
rect 21088 26732 21140 26741
rect 27620 26868 27672 26920
rect 29000 26936 29052 26988
rect 29920 27004 29972 27056
rect 29552 26979 29604 26988
rect 29552 26945 29561 26979
rect 29561 26945 29595 26979
rect 29595 26945 29604 26979
rect 29552 26936 29604 26945
rect 30012 26936 30064 26988
rect 30196 26936 30248 26988
rect 31300 27004 31352 27056
rect 32864 27004 32916 27056
rect 33600 26936 33652 26988
rect 36820 27004 36872 27056
rect 35348 26936 35400 26988
rect 36360 26979 36412 26988
rect 36360 26945 36369 26979
rect 36369 26945 36403 26979
rect 36403 26945 36412 26979
rect 36360 26936 36412 26945
rect 36452 26979 36504 26988
rect 36452 26945 36461 26979
rect 36461 26945 36495 26979
rect 36495 26945 36504 26979
rect 36636 26979 36688 26988
rect 36452 26936 36504 26945
rect 36636 26945 36645 26979
rect 36645 26945 36679 26979
rect 36679 26945 36688 26979
rect 36636 26936 36688 26945
rect 37556 27072 37608 27124
rect 37648 26979 37700 26988
rect 37648 26945 37657 26979
rect 37657 26945 37691 26979
rect 37691 26945 37700 26979
rect 37648 26936 37700 26945
rect 24676 26732 24728 26784
rect 26424 26732 26476 26784
rect 26516 26775 26568 26784
rect 26516 26741 26525 26775
rect 26525 26741 26559 26775
rect 26559 26741 26568 26775
rect 26516 26732 26568 26741
rect 30104 26732 30156 26784
rect 38016 26868 38068 26920
rect 36912 26800 36964 26852
rect 35532 26732 35584 26784
rect 36176 26775 36228 26784
rect 36176 26741 36185 26775
rect 36185 26741 36219 26775
rect 36219 26741 36228 26775
rect 36176 26732 36228 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18328 26528 18380 26580
rect 19064 26528 19116 26580
rect 21364 26571 21416 26580
rect 21364 26537 21373 26571
rect 21373 26537 21407 26571
rect 21407 26537 21416 26571
rect 21364 26528 21416 26537
rect 26148 26528 26200 26580
rect 27712 26528 27764 26580
rect 27896 26528 27948 26580
rect 29000 26571 29052 26580
rect 29000 26537 29009 26571
rect 29009 26537 29043 26571
rect 29043 26537 29052 26571
rect 29000 26528 29052 26537
rect 36360 26528 36412 26580
rect 33324 26460 33376 26512
rect 34612 26460 34664 26512
rect 18236 26392 18288 26444
rect 18788 26435 18840 26444
rect 18788 26401 18797 26435
rect 18797 26401 18831 26435
rect 18831 26401 18840 26435
rect 18788 26392 18840 26401
rect 30380 26435 30432 26444
rect 30380 26401 30389 26435
rect 30389 26401 30423 26435
rect 30423 26401 30432 26435
rect 30380 26392 30432 26401
rect 32588 26392 32640 26444
rect 17960 26324 18012 26376
rect 18512 26367 18564 26376
rect 17224 26256 17276 26308
rect 17776 26256 17828 26308
rect 18512 26333 18521 26367
rect 18521 26333 18555 26367
rect 18555 26333 18564 26367
rect 18512 26324 18564 26333
rect 21088 26324 21140 26376
rect 23112 26367 23164 26376
rect 19248 26256 19300 26308
rect 20076 26256 20128 26308
rect 23112 26333 23121 26367
rect 23121 26333 23155 26367
rect 23155 26333 23164 26367
rect 23112 26324 23164 26333
rect 24676 26324 24728 26376
rect 26240 26324 26292 26376
rect 27160 26324 27212 26376
rect 28540 26324 28592 26376
rect 29000 26324 29052 26376
rect 30104 26367 30156 26376
rect 30104 26333 30113 26367
rect 30113 26333 30147 26367
rect 30147 26333 30156 26367
rect 30104 26324 30156 26333
rect 30288 26367 30340 26376
rect 30288 26333 30297 26367
rect 30297 26333 30331 26367
rect 30331 26333 30340 26367
rect 30288 26324 30340 26333
rect 33600 26367 33652 26376
rect 33600 26333 33609 26367
rect 33609 26333 33643 26367
rect 33643 26333 33652 26367
rect 33600 26324 33652 26333
rect 35348 26392 35400 26444
rect 36176 26392 36228 26444
rect 36820 26392 36872 26444
rect 35256 26367 35308 26376
rect 35256 26333 35265 26367
rect 35265 26333 35299 26367
rect 35299 26333 35308 26367
rect 35256 26324 35308 26333
rect 35624 26324 35676 26376
rect 24492 26256 24544 26308
rect 25596 26256 25648 26308
rect 30196 26256 30248 26308
rect 31208 26299 31260 26308
rect 31208 26265 31217 26299
rect 31217 26265 31251 26299
rect 31251 26265 31260 26299
rect 31208 26256 31260 26265
rect 33692 26256 33744 26308
rect 34612 26256 34664 26308
rect 35808 26256 35860 26308
rect 36176 26256 36228 26308
rect 22928 26188 22980 26240
rect 32036 26188 32088 26240
rect 34888 26231 34940 26240
rect 34888 26197 34897 26231
rect 34897 26197 34931 26231
rect 34931 26197 34940 26231
rect 34888 26188 34940 26197
rect 37280 26188 37332 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 23112 25984 23164 26036
rect 24676 26027 24728 26036
rect 24676 25993 24685 26027
rect 24685 25993 24719 26027
rect 24719 25993 24728 26027
rect 24676 25984 24728 25993
rect 25596 26027 25648 26036
rect 25596 25993 25605 26027
rect 25605 25993 25639 26027
rect 25639 25993 25648 26027
rect 25596 25984 25648 25993
rect 29644 25984 29696 26036
rect 19340 25916 19392 25968
rect 16948 25848 17000 25900
rect 19708 25891 19760 25900
rect 19708 25857 19717 25891
rect 19717 25857 19751 25891
rect 19751 25857 19760 25891
rect 19708 25848 19760 25857
rect 22192 25916 22244 25968
rect 22560 25959 22612 25968
rect 22560 25925 22569 25959
rect 22569 25925 22603 25959
rect 22603 25925 22612 25959
rect 22560 25916 22612 25925
rect 20076 25891 20128 25900
rect 17500 25823 17552 25832
rect 17500 25789 17509 25823
rect 17509 25789 17543 25823
rect 17543 25789 17552 25823
rect 17500 25780 17552 25789
rect 19340 25780 19392 25832
rect 20076 25857 20085 25891
rect 20085 25857 20119 25891
rect 20119 25857 20128 25891
rect 20076 25848 20128 25857
rect 23112 25848 23164 25900
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 26516 25916 26568 25968
rect 30196 25916 30248 25968
rect 34428 25984 34480 26036
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 28816 25848 28868 25900
rect 31392 25848 31444 25900
rect 34520 25916 34572 25968
rect 34796 25916 34848 25968
rect 35256 25916 35308 25968
rect 34888 25848 34940 25900
rect 24400 25780 24452 25832
rect 24952 25780 25004 25832
rect 26332 25780 26384 25832
rect 29368 25823 29420 25832
rect 29368 25789 29377 25823
rect 29377 25789 29411 25823
rect 29411 25789 29420 25823
rect 29368 25780 29420 25789
rect 29828 25823 29880 25832
rect 29828 25789 29837 25823
rect 29837 25789 29871 25823
rect 29871 25789 29880 25823
rect 29828 25780 29880 25789
rect 34796 25823 34848 25832
rect 34796 25789 34805 25823
rect 34805 25789 34839 25823
rect 34839 25789 34848 25823
rect 34796 25780 34848 25789
rect 17960 25755 18012 25764
rect 17960 25721 17969 25755
rect 17969 25721 18003 25755
rect 18003 25721 18012 25755
rect 17960 25712 18012 25721
rect 31024 25712 31076 25764
rect 36176 25984 36228 26036
rect 37464 25984 37516 26036
rect 37648 25891 37700 25900
rect 37648 25857 37657 25891
rect 37657 25857 37691 25891
rect 37691 25857 37700 25891
rect 37648 25848 37700 25857
rect 36636 25780 36688 25832
rect 37188 25780 37240 25832
rect 20076 25644 20128 25696
rect 23204 25644 23256 25696
rect 29184 25687 29236 25696
rect 29184 25653 29193 25687
rect 29193 25653 29227 25687
rect 29227 25653 29236 25687
rect 29184 25644 29236 25653
rect 30748 25644 30800 25696
rect 35348 25644 35400 25696
rect 37004 25644 37056 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 17224 25483 17276 25492
rect 17224 25449 17233 25483
rect 17233 25449 17267 25483
rect 17267 25449 17276 25483
rect 17224 25440 17276 25449
rect 19708 25440 19760 25492
rect 22100 25440 22152 25492
rect 22560 25440 22612 25492
rect 22468 25372 22520 25424
rect 17316 25304 17368 25356
rect 17960 25304 18012 25356
rect 19064 25304 19116 25356
rect 17408 25279 17460 25288
rect 17408 25245 17417 25279
rect 17417 25245 17451 25279
rect 17451 25245 17460 25279
rect 17408 25236 17460 25245
rect 17684 25279 17736 25288
rect 17684 25245 17693 25279
rect 17693 25245 17727 25279
rect 17727 25245 17736 25279
rect 18236 25279 18288 25288
rect 17684 25236 17736 25245
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 18788 25236 18840 25288
rect 19892 25236 19944 25288
rect 20076 25279 20128 25288
rect 20076 25245 20110 25279
rect 20110 25245 20128 25279
rect 20076 25236 20128 25245
rect 21916 25304 21968 25356
rect 24492 25440 24544 25492
rect 27160 25483 27212 25492
rect 27160 25449 27169 25483
rect 27169 25449 27203 25483
rect 27203 25449 27212 25483
rect 27160 25440 27212 25449
rect 29000 25483 29052 25492
rect 29000 25449 29009 25483
rect 29009 25449 29043 25483
rect 29043 25449 29052 25483
rect 29000 25440 29052 25449
rect 29276 25440 29328 25492
rect 29368 25440 29420 25492
rect 31392 25483 31444 25492
rect 24584 25372 24636 25424
rect 21824 25279 21876 25288
rect 21824 25245 21833 25279
rect 21833 25245 21867 25279
rect 21867 25245 21876 25279
rect 21824 25236 21876 25245
rect 22652 25279 22704 25288
rect 22652 25245 22661 25279
rect 22661 25245 22695 25279
rect 22695 25245 22704 25279
rect 22652 25236 22704 25245
rect 22928 25279 22980 25288
rect 22928 25245 22962 25279
rect 22962 25245 22980 25279
rect 22928 25236 22980 25245
rect 23204 25236 23256 25288
rect 24492 25236 24544 25288
rect 24860 25347 24912 25356
rect 24860 25313 24869 25347
rect 24869 25313 24903 25347
rect 24903 25313 24912 25347
rect 26332 25372 26384 25424
rect 24860 25304 24912 25313
rect 26240 25304 26292 25356
rect 31392 25449 31401 25483
rect 31401 25449 31435 25483
rect 31435 25449 31444 25483
rect 31392 25440 31444 25449
rect 33324 25440 33376 25492
rect 33508 25440 33560 25492
rect 34060 25483 34112 25492
rect 34060 25449 34069 25483
rect 34069 25449 34103 25483
rect 34103 25449 34112 25483
rect 34060 25440 34112 25449
rect 19248 25168 19300 25220
rect 21364 25168 21416 25220
rect 23112 25168 23164 25220
rect 24768 25168 24820 25220
rect 25872 25236 25924 25288
rect 26516 25236 26568 25288
rect 27804 25279 27856 25288
rect 27804 25245 27813 25279
rect 27813 25245 27847 25279
rect 27847 25245 27856 25279
rect 27804 25236 27856 25245
rect 29000 25304 29052 25356
rect 29828 25304 29880 25356
rect 36728 25304 36780 25356
rect 18604 25100 18656 25152
rect 22008 25100 22060 25152
rect 22284 25100 22336 25152
rect 26516 25143 26568 25152
rect 26516 25109 26525 25143
rect 26525 25109 26559 25143
rect 26559 25109 26568 25143
rect 26516 25100 26568 25109
rect 27620 25168 27672 25220
rect 27896 25143 27948 25152
rect 27896 25109 27905 25143
rect 27905 25109 27939 25143
rect 27939 25109 27948 25143
rect 27896 25100 27948 25109
rect 28816 25211 28868 25220
rect 28816 25177 28825 25211
rect 28825 25177 28859 25211
rect 28859 25177 28868 25211
rect 28816 25168 28868 25177
rect 29368 25168 29420 25220
rect 30840 25168 30892 25220
rect 32956 25168 33008 25220
rect 33324 25168 33376 25220
rect 34520 25236 34572 25288
rect 36176 25236 36228 25288
rect 37004 25236 37056 25288
rect 34980 25168 35032 25220
rect 30012 25100 30064 25152
rect 33876 25100 33928 25152
rect 37188 25100 37240 25152
rect 37648 25100 37700 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 16304 24803 16356 24812
rect 16304 24769 16313 24803
rect 16313 24769 16347 24803
rect 16347 24769 16356 24803
rect 17408 24828 17460 24880
rect 17868 24828 17920 24880
rect 16304 24760 16356 24769
rect 17776 24803 17828 24812
rect 17776 24769 17785 24803
rect 17785 24769 17819 24803
rect 17819 24769 17828 24803
rect 17776 24760 17828 24769
rect 22008 24896 22060 24948
rect 24492 24896 24544 24948
rect 27620 24896 27672 24948
rect 28540 24939 28592 24948
rect 28540 24905 28549 24939
rect 28549 24905 28583 24939
rect 28583 24905 28592 24939
rect 28540 24896 28592 24905
rect 34980 24896 35032 24948
rect 37188 24896 37240 24948
rect 18604 24803 18656 24812
rect 18604 24769 18613 24803
rect 18613 24769 18647 24803
rect 18647 24769 18656 24803
rect 18604 24760 18656 24769
rect 18788 24760 18840 24812
rect 19064 24803 19116 24812
rect 19064 24769 19073 24803
rect 19073 24769 19107 24803
rect 19107 24769 19116 24803
rect 19064 24760 19116 24769
rect 18696 24692 18748 24744
rect 17040 24624 17092 24676
rect 19984 24760 20036 24812
rect 20168 24803 20220 24812
rect 20168 24769 20202 24803
rect 20202 24769 20220 24803
rect 20168 24760 20220 24769
rect 22100 24760 22152 24812
rect 22468 24760 22520 24812
rect 24676 24828 24728 24880
rect 24492 24760 24544 24812
rect 26516 24828 26568 24880
rect 19340 24624 19392 24676
rect 17316 24556 17368 24608
rect 18788 24556 18840 24608
rect 21824 24692 21876 24744
rect 22652 24624 22704 24676
rect 25964 24803 26016 24812
rect 25964 24769 25973 24803
rect 25973 24769 26007 24803
rect 26007 24769 26016 24803
rect 25964 24760 26016 24769
rect 26424 24760 26476 24812
rect 27896 24760 27948 24812
rect 28540 24760 28592 24812
rect 30748 24760 30800 24812
rect 26332 24692 26384 24744
rect 29000 24735 29052 24744
rect 29000 24701 29009 24735
rect 29009 24701 29043 24735
rect 29043 24701 29052 24735
rect 29000 24692 29052 24701
rect 30012 24692 30064 24744
rect 30288 24692 30340 24744
rect 32312 24760 32364 24812
rect 33876 24828 33928 24880
rect 33692 24803 33744 24812
rect 31944 24692 31996 24744
rect 33692 24769 33701 24803
rect 33701 24769 33735 24803
rect 33735 24769 33744 24803
rect 33692 24760 33744 24769
rect 35348 24760 35400 24812
rect 38292 24828 38344 24880
rect 37464 24803 37516 24812
rect 37464 24769 37473 24803
rect 37473 24769 37507 24803
rect 37507 24769 37516 24803
rect 37464 24760 37516 24769
rect 37648 24760 37700 24812
rect 33416 24692 33468 24744
rect 37556 24692 37608 24744
rect 30840 24667 30892 24676
rect 30840 24633 30849 24667
rect 30849 24633 30883 24667
rect 30883 24633 30892 24667
rect 30840 24624 30892 24633
rect 32956 24624 33008 24676
rect 36912 24667 36964 24676
rect 36912 24633 36921 24667
rect 36921 24633 36955 24667
rect 36955 24633 36964 24667
rect 36912 24624 36964 24633
rect 37280 24624 37332 24676
rect 21272 24599 21324 24608
rect 21272 24565 21281 24599
rect 21281 24565 21315 24599
rect 21315 24565 21324 24599
rect 21272 24556 21324 24565
rect 25412 24556 25464 24608
rect 25872 24556 25924 24608
rect 29276 24556 29328 24608
rect 32128 24556 32180 24608
rect 32588 24599 32640 24608
rect 32588 24565 32597 24599
rect 32597 24565 32631 24599
rect 32631 24565 32640 24599
rect 32588 24556 32640 24565
rect 33048 24599 33100 24608
rect 33048 24565 33057 24599
rect 33057 24565 33091 24599
rect 33091 24565 33100 24599
rect 33048 24556 33100 24565
rect 37188 24556 37240 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 16304 24352 16356 24404
rect 16948 24191 17000 24200
rect 16948 24157 16957 24191
rect 16957 24157 16991 24191
rect 16991 24157 17000 24191
rect 16948 24148 17000 24157
rect 17684 24352 17736 24404
rect 20168 24352 20220 24404
rect 22284 24395 22336 24404
rect 22284 24361 22293 24395
rect 22293 24361 22327 24395
rect 22327 24361 22336 24395
rect 22284 24352 22336 24361
rect 24492 24352 24544 24404
rect 26240 24352 26292 24404
rect 26516 24352 26568 24404
rect 27804 24352 27856 24404
rect 28540 24395 28592 24404
rect 28540 24361 28549 24395
rect 28549 24361 28583 24395
rect 28583 24361 28592 24395
rect 28540 24352 28592 24361
rect 17316 24284 17368 24336
rect 17224 24259 17276 24268
rect 17224 24225 17233 24259
rect 17233 24225 17267 24259
rect 17267 24225 17276 24259
rect 17224 24216 17276 24225
rect 17500 24216 17552 24268
rect 23756 24327 23808 24336
rect 23756 24293 23765 24327
rect 23765 24293 23799 24327
rect 23799 24293 23808 24327
rect 23756 24284 23808 24293
rect 29184 24352 29236 24404
rect 33416 24395 33468 24404
rect 33416 24361 33425 24395
rect 33425 24361 33459 24395
rect 33459 24361 33468 24395
rect 33416 24352 33468 24361
rect 37556 24395 37608 24404
rect 37556 24361 37565 24395
rect 37565 24361 37599 24395
rect 37599 24361 37608 24395
rect 37556 24352 37608 24361
rect 29368 24284 29420 24336
rect 19432 24216 19484 24268
rect 17868 24191 17920 24200
rect 17868 24157 17877 24191
rect 17877 24157 17911 24191
rect 17911 24157 17920 24191
rect 17868 24148 17920 24157
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 18788 24148 18840 24200
rect 19984 24191 20036 24200
rect 19984 24157 19993 24191
rect 19993 24157 20027 24191
rect 20027 24157 20036 24191
rect 19984 24148 20036 24157
rect 20260 24148 20312 24200
rect 21272 24148 21324 24200
rect 21640 24191 21692 24200
rect 21640 24157 21649 24191
rect 21649 24157 21683 24191
rect 21683 24157 21692 24191
rect 21640 24148 21692 24157
rect 22560 24216 22612 24268
rect 22008 24191 22060 24200
rect 22008 24157 22017 24191
rect 22017 24157 22051 24191
rect 22051 24157 22060 24191
rect 22008 24148 22060 24157
rect 22100 24148 22152 24200
rect 23204 24216 23256 24268
rect 23572 24216 23624 24268
rect 23112 24191 23164 24200
rect 23112 24157 23121 24191
rect 23121 24157 23155 24191
rect 23155 24157 23164 24191
rect 23112 24148 23164 24157
rect 24676 24216 24728 24268
rect 26332 24216 26384 24268
rect 18236 24055 18288 24064
rect 18236 24021 18245 24055
rect 18245 24021 18279 24055
rect 18279 24021 18288 24055
rect 18236 24012 18288 24021
rect 23848 24080 23900 24132
rect 24584 24191 24636 24200
rect 24584 24157 24593 24191
rect 24593 24157 24627 24191
rect 24627 24157 24636 24191
rect 24584 24148 24636 24157
rect 24768 24191 24820 24200
rect 24768 24157 24777 24191
rect 24777 24157 24811 24191
rect 24811 24157 24820 24191
rect 24768 24148 24820 24157
rect 25412 24148 25464 24200
rect 27620 24148 27672 24200
rect 28724 24191 28776 24200
rect 28724 24157 28733 24191
rect 28733 24157 28767 24191
rect 28767 24157 28776 24191
rect 28724 24148 28776 24157
rect 29276 24148 29328 24200
rect 31760 24216 31812 24268
rect 36176 24259 36228 24268
rect 36176 24225 36185 24259
rect 36185 24225 36219 24259
rect 36219 24225 36228 24259
rect 36176 24216 36228 24225
rect 32036 24191 32088 24200
rect 32036 24157 32045 24191
rect 32045 24157 32079 24191
rect 32079 24157 32088 24191
rect 32036 24148 32088 24157
rect 32128 24148 32180 24200
rect 33876 24080 33928 24132
rect 22376 24012 22428 24064
rect 22468 24012 22520 24064
rect 31392 24055 31444 24064
rect 31392 24021 31401 24055
rect 31401 24021 31435 24055
rect 31435 24021 31444 24055
rect 31392 24012 31444 24021
rect 31760 24012 31812 24064
rect 36636 24080 36688 24132
rect 34796 24012 34848 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 17224 23808 17276 23860
rect 19984 23808 20036 23860
rect 21640 23808 21692 23860
rect 28724 23808 28776 23860
rect 29184 23808 29236 23860
rect 32864 23808 32916 23860
rect 36636 23851 36688 23860
rect 17776 23740 17828 23792
rect 23388 23783 23440 23792
rect 18236 23672 18288 23724
rect 19432 23715 19484 23724
rect 19432 23681 19441 23715
rect 19441 23681 19475 23715
rect 19475 23681 19484 23715
rect 19432 23672 19484 23681
rect 21272 23715 21324 23724
rect 21272 23681 21281 23715
rect 21281 23681 21315 23715
rect 21315 23681 21324 23715
rect 21272 23672 21324 23681
rect 23388 23749 23397 23783
rect 23397 23749 23431 23783
rect 23431 23749 23440 23783
rect 23388 23740 23440 23749
rect 22008 23715 22060 23724
rect 22008 23681 22017 23715
rect 22017 23681 22051 23715
rect 22051 23681 22060 23715
rect 22008 23672 22060 23681
rect 22192 23715 22244 23724
rect 22192 23681 22201 23715
rect 22201 23681 22235 23715
rect 22235 23681 22244 23715
rect 22192 23672 22244 23681
rect 22376 23715 22428 23724
rect 22376 23681 22385 23715
rect 22385 23681 22419 23715
rect 22419 23681 22428 23715
rect 22376 23672 22428 23681
rect 22560 23715 22612 23724
rect 22560 23681 22569 23715
rect 22569 23681 22603 23715
rect 22603 23681 22612 23715
rect 22560 23672 22612 23681
rect 25964 23715 26016 23724
rect 25964 23681 25973 23715
rect 25973 23681 26007 23715
rect 26007 23681 26016 23715
rect 25964 23672 26016 23681
rect 26240 23672 26292 23724
rect 26976 23672 27028 23724
rect 31392 23740 31444 23792
rect 29460 23672 29512 23724
rect 21824 23604 21876 23656
rect 29092 23604 29144 23656
rect 32036 23672 32088 23724
rect 32956 23740 33008 23792
rect 36636 23817 36645 23851
rect 36645 23817 36679 23851
rect 36679 23817 36688 23851
rect 36636 23808 36688 23817
rect 35532 23783 35584 23792
rect 35532 23749 35541 23783
rect 35541 23749 35575 23783
rect 35575 23749 35584 23783
rect 35532 23740 35584 23749
rect 36176 23740 36228 23792
rect 33784 23715 33836 23724
rect 33784 23681 33793 23715
rect 33793 23681 33827 23715
rect 33827 23681 33836 23715
rect 33784 23672 33836 23681
rect 37280 23672 37332 23724
rect 37464 23715 37516 23724
rect 37464 23681 37473 23715
rect 37473 23681 37507 23715
rect 37507 23681 37516 23715
rect 37464 23672 37516 23681
rect 37648 23715 37700 23724
rect 37648 23681 37657 23715
rect 37657 23681 37691 23715
rect 37691 23681 37700 23715
rect 37648 23672 37700 23681
rect 22652 23536 22704 23588
rect 33416 23604 33468 23656
rect 34244 23536 34296 23588
rect 21640 23468 21692 23520
rect 26240 23511 26292 23520
rect 26240 23477 26249 23511
rect 26249 23477 26283 23511
rect 26283 23477 26292 23511
rect 26240 23468 26292 23477
rect 31944 23468 31996 23520
rect 32588 23511 32640 23520
rect 32588 23477 32597 23511
rect 32597 23477 32631 23511
rect 32631 23477 32640 23511
rect 32588 23468 32640 23477
rect 37556 23468 37608 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 19432 23264 19484 23316
rect 20444 23264 20496 23316
rect 22008 23264 22060 23316
rect 23848 23264 23900 23316
rect 20812 23171 20864 23180
rect 20812 23137 20821 23171
rect 20821 23137 20855 23171
rect 20855 23137 20864 23171
rect 20812 23128 20864 23137
rect 22652 23171 22704 23180
rect 22652 23137 22661 23171
rect 22661 23137 22695 23171
rect 22695 23137 22704 23171
rect 22652 23128 22704 23137
rect 17776 23103 17828 23112
rect 17776 23069 17785 23103
rect 17785 23069 17819 23103
rect 17819 23069 17828 23103
rect 17776 23060 17828 23069
rect 18604 23035 18656 23044
rect 18604 23001 18613 23035
rect 18613 23001 18647 23035
rect 18647 23001 18656 23035
rect 19340 23060 19392 23112
rect 19984 23060 20036 23112
rect 20720 23103 20772 23112
rect 20720 23069 20729 23103
rect 20729 23069 20763 23103
rect 20763 23069 20772 23103
rect 20720 23060 20772 23069
rect 18604 22992 18656 23001
rect 21272 22992 21324 23044
rect 21640 23103 21692 23112
rect 21640 23069 21649 23103
rect 21649 23069 21683 23103
rect 21683 23069 21692 23103
rect 21824 23103 21876 23112
rect 21640 23060 21692 23069
rect 21824 23069 21833 23103
rect 21833 23069 21867 23103
rect 21867 23069 21876 23103
rect 21824 23060 21876 23069
rect 21916 23103 21968 23112
rect 21916 23069 21935 23103
rect 21935 23069 21968 23103
rect 21916 23060 21968 23069
rect 22192 22992 22244 23044
rect 22928 23035 22980 23044
rect 22928 23001 22962 23035
rect 22962 23001 22980 23035
rect 22928 22992 22980 23001
rect 17960 22967 18012 22976
rect 17960 22933 17969 22967
rect 17969 22933 18003 22967
rect 18003 22933 18012 22967
rect 17960 22924 18012 22933
rect 18788 22967 18840 22976
rect 18788 22933 18797 22967
rect 18797 22933 18831 22967
rect 18831 22933 18840 22967
rect 18788 22924 18840 22933
rect 19340 22924 19392 22976
rect 20260 22924 20312 22976
rect 21364 22924 21416 22976
rect 31208 23307 31260 23316
rect 31208 23273 31217 23307
rect 31217 23273 31251 23307
rect 31251 23273 31260 23307
rect 31208 23264 31260 23273
rect 33784 23264 33836 23316
rect 34244 23307 34296 23316
rect 32312 23239 32364 23248
rect 26240 23128 26292 23180
rect 26332 23171 26384 23180
rect 26332 23137 26341 23171
rect 26341 23137 26375 23171
rect 26375 23137 26384 23171
rect 26332 23128 26384 23137
rect 25964 22992 26016 23044
rect 26792 23060 26844 23112
rect 32312 23205 32321 23239
rect 32321 23205 32355 23239
rect 32355 23205 32364 23239
rect 32312 23196 32364 23205
rect 32864 23196 32916 23248
rect 31944 23171 31996 23180
rect 31944 23137 31953 23171
rect 31953 23137 31987 23171
rect 31987 23137 31996 23171
rect 34244 23273 34253 23307
rect 34253 23273 34287 23307
rect 34287 23273 34296 23307
rect 34244 23264 34296 23273
rect 38292 23307 38344 23316
rect 38292 23273 38301 23307
rect 38301 23273 38335 23307
rect 38335 23273 38344 23307
rect 38292 23264 38344 23273
rect 31944 23128 31996 23137
rect 36176 23128 36228 23180
rect 25688 22924 25740 22976
rect 29000 23060 29052 23112
rect 31760 23060 31812 23112
rect 33048 23103 33100 23112
rect 33048 23069 33057 23103
rect 33057 23069 33091 23103
rect 33091 23069 33100 23103
rect 33048 23060 33100 23069
rect 29092 22992 29144 23044
rect 33140 23069 33149 23078
rect 33149 23069 33183 23078
rect 33183 23069 33192 23078
rect 33140 23026 33192 23069
rect 33508 23060 33560 23112
rect 34888 23103 34940 23112
rect 34888 23069 34897 23103
rect 34897 23069 34931 23103
rect 34931 23069 34940 23103
rect 34888 23060 34940 23069
rect 35532 23060 35584 23112
rect 33692 22992 33744 23044
rect 33876 23035 33928 23044
rect 33876 23001 33885 23035
rect 33885 23001 33919 23035
rect 33919 23001 33928 23035
rect 33876 22992 33928 23001
rect 34520 22992 34572 23044
rect 34796 22992 34848 23044
rect 37372 22992 37424 23044
rect 35532 22924 35584 22976
rect 35808 22924 35860 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 17868 22763 17920 22772
rect 17868 22729 17877 22763
rect 17877 22729 17911 22763
rect 17911 22729 17920 22763
rect 17868 22720 17920 22729
rect 18052 22720 18104 22772
rect 17960 22584 18012 22636
rect 18144 22584 18196 22636
rect 18788 22720 18840 22772
rect 19432 22720 19484 22772
rect 21272 22720 21324 22772
rect 21824 22720 21876 22772
rect 18604 22584 18656 22636
rect 19156 22627 19208 22636
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 19064 22516 19116 22568
rect 22376 22652 22428 22704
rect 22928 22720 22980 22772
rect 25688 22763 25740 22772
rect 25688 22729 25697 22763
rect 25697 22729 25731 22763
rect 25731 22729 25740 22763
rect 25688 22720 25740 22729
rect 26332 22720 26384 22772
rect 30564 22763 30616 22772
rect 30564 22729 30573 22763
rect 30573 22729 30607 22763
rect 30607 22729 30616 22763
rect 30564 22720 30616 22729
rect 33692 22763 33744 22772
rect 33692 22729 33701 22763
rect 33701 22729 33735 22763
rect 33735 22729 33744 22763
rect 33692 22720 33744 22729
rect 33968 22720 34020 22772
rect 23572 22652 23624 22704
rect 24032 22652 24084 22704
rect 24400 22652 24452 22704
rect 23112 22584 23164 22636
rect 23756 22584 23808 22636
rect 24584 22627 24636 22636
rect 24584 22593 24618 22627
rect 24618 22593 24636 22627
rect 24584 22584 24636 22593
rect 27988 22627 28040 22636
rect 27988 22593 28022 22627
rect 28022 22593 28040 22627
rect 31116 22652 31168 22704
rect 32588 22695 32640 22704
rect 32588 22661 32622 22695
rect 32622 22661 32640 22695
rect 32588 22652 32640 22661
rect 37280 22720 37332 22772
rect 27988 22584 28040 22593
rect 30288 22627 30340 22636
rect 30288 22593 30297 22627
rect 30297 22593 30331 22627
rect 30331 22593 30340 22627
rect 30288 22584 30340 22593
rect 19432 22516 19484 22568
rect 24308 22559 24360 22568
rect 24308 22525 24317 22559
rect 24317 22525 24351 22559
rect 24351 22525 24360 22559
rect 24308 22516 24360 22525
rect 25780 22516 25832 22568
rect 23112 22448 23164 22500
rect 26516 22516 26568 22568
rect 27712 22559 27764 22568
rect 19984 22380 20036 22432
rect 21364 22380 21416 22432
rect 22192 22380 22244 22432
rect 22560 22380 22612 22432
rect 27712 22525 27721 22559
rect 27721 22525 27755 22559
rect 27755 22525 27764 22559
rect 27712 22516 27764 22525
rect 30564 22448 30616 22500
rect 31484 22423 31536 22432
rect 31484 22389 31493 22423
rect 31493 22389 31527 22423
rect 31527 22389 31536 22423
rect 31484 22380 31536 22389
rect 32036 22584 32088 22636
rect 33140 22584 33192 22636
rect 34428 22627 34480 22636
rect 33416 22380 33468 22432
rect 34428 22593 34437 22627
rect 34437 22593 34471 22627
rect 34471 22593 34480 22627
rect 34428 22584 34480 22593
rect 34888 22627 34940 22636
rect 34888 22593 34897 22627
rect 34897 22593 34931 22627
rect 34931 22593 34940 22627
rect 34888 22584 34940 22593
rect 38292 22652 38344 22704
rect 37648 22627 37700 22636
rect 37648 22593 37657 22627
rect 37657 22593 37691 22627
rect 37691 22593 37700 22627
rect 37648 22584 37700 22593
rect 35624 22380 35676 22432
rect 36268 22423 36320 22432
rect 36268 22389 36277 22423
rect 36277 22389 36311 22423
rect 36311 22389 36320 22423
rect 36268 22380 36320 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 18788 22176 18840 22228
rect 20444 22219 20496 22228
rect 20444 22185 20453 22219
rect 20453 22185 20487 22219
rect 20487 22185 20496 22219
rect 20444 22176 20496 22185
rect 17868 22040 17920 22092
rect 17960 22015 18012 22024
rect 17960 21981 17969 22015
rect 17969 21981 18003 22015
rect 18003 21981 18012 22015
rect 17960 21972 18012 21981
rect 18144 21904 18196 21956
rect 20720 21972 20772 22024
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 21364 21972 21416 22024
rect 22560 22015 22612 22024
rect 22560 21981 22569 22015
rect 22569 21981 22603 22015
rect 22603 21981 22612 22015
rect 22560 21972 22612 21981
rect 23112 21972 23164 22024
rect 24584 22176 24636 22228
rect 23572 21972 23624 22024
rect 26516 22083 26568 22092
rect 26516 22049 26525 22083
rect 26525 22049 26559 22083
rect 26559 22049 26568 22083
rect 26516 22040 26568 22049
rect 25780 22015 25832 22024
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21972 25832 21981
rect 26792 21972 26844 22024
rect 18052 21836 18104 21888
rect 20904 21904 20956 21956
rect 25228 21904 25280 21956
rect 26976 22151 27028 22160
rect 26976 22117 26985 22151
rect 26985 22117 27019 22151
rect 27019 22117 27028 22151
rect 26976 22108 27028 22117
rect 18880 21836 18932 21888
rect 20076 21879 20128 21888
rect 20076 21845 20085 21879
rect 20085 21845 20119 21879
rect 20119 21845 20128 21879
rect 20076 21836 20128 21845
rect 22100 21879 22152 21888
rect 22100 21845 22109 21879
rect 22109 21845 22143 21879
rect 22143 21845 22152 21879
rect 23204 21879 23256 21888
rect 22100 21836 22152 21845
rect 23204 21845 23213 21879
rect 23213 21845 23247 21879
rect 23247 21845 23256 21879
rect 23204 21836 23256 21845
rect 29092 22176 29144 22228
rect 31760 22176 31812 22228
rect 28540 22015 28592 22024
rect 28540 21981 28549 22015
rect 28549 21981 28583 22015
rect 28583 21981 28592 22015
rect 28540 21972 28592 21981
rect 33140 22040 33192 22092
rect 34428 22176 34480 22228
rect 35164 22176 35216 22228
rect 35808 22176 35860 22228
rect 37372 22219 37424 22228
rect 37372 22185 37381 22219
rect 37381 22185 37415 22219
rect 37415 22185 37424 22219
rect 37372 22176 37424 22185
rect 34704 22040 34756 22092
rect 35532 22083 35584 22092
rect 35532 22049 35541 22083
rect 35541 22049 35575 22083
rect 35575 22049 35584 22083
rect 35532 22040 35584 22049
rect 36176 22083 36228 22092
rect 29000 21972 29052 22024
rect 30012 22015 30064 22024
rect 30012 21981 30021 22015
rect 30021 21981 30055 22015
rect 30055 21981 30064 22015
rect 30012 21972 30064 21981
rect 31484 21972 31536 22024
rect 32496 22015 32548 22024
rect 32496 21981 32505 22015
rect 32505 21981 32539 22015
rect 32539 21981 32548 22015
rect 32496 21972 32548 21981
rect 32588 22015 32640 22024
rect 32588 21981 32597 22015
rect 32597 21981 32631 22015
rect 32631 21981 32640 22015
rect 32588 21972 32640 21981
rect 33600 21972 33652 22024
rect 31392 21879 31444 21888
rect 31392 21845 31401 21879
rect 31401 21845 31435 21879
rect 31435 21845 31444 21879
rect 31392 21836 31444 21845
rect 33508 21904 33560 21956
rect 34152 22015 34204 22024
rect 34152 21981 34161 22015
rect 34161 21981 34195 22015
rect 34195 21981 34204 22015
rect 34152 21972 34204 21981
rect 35900 21972 35952 22024
rect 36176 22049 36185 22083
rect 36185 22049 36219 22083
rect 36219 22049 36228 22083
rect 36176 22040 36228 22049
rect 36268 22015 36320 22024
rect 36268 21981 36277 22015
rect 36277 21981 36311 22015
rect 36311 21981 36320 22015
rect 36268 21972 36320 21981
rect 37556 22015 37608 22024
rect 37556 21981 37565 22015
rect 37565 21981 37599 22015
rect 37599 21981 37608 22015
rect 37556 21972 37608 21981
rect 35164 21947 35216 21956
rect 35164 21913 35173 21947
rect 35173 21913 35207 21947
rect 35207 21913 35216 21947
rect 35164 21904 35216 21913
rect 35348 21879 35400 21888
rect 35348 21845 35357 21879
rect 35357 21845 35391 21879
rect 35391 21845 35400 21879
rect 35348 21836 35400 21845
rect 35624 21836 35676 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 19064 21632 19116 21684
rect 21180 21675 21232 21684
rect 21180 21641 21189 21675
rect 21189 21641 21223 21675
rect 21223 21641 21232 21675
rect 21180 21632 21232 21641
rect 23204 21632 23256 21684
rect 27988 21675 28040 21684
rect 27988 21641 27997 21675
rect 27997 21641 28031 21675
rect 28031 21641 28040 21675
rect 27988 21632 28040 21641
rect 28540 21632 28592 21684
rect 17868 21496 17920 21548
rect 18788 21496 18840 21548
rect 19432 21496 19484 21548
rect 22100 21564 22152 21616
rect 19892 21496 19944 21548
rect 20076 21539 20128 21548
rect 20076 21505 20110 21539
rect 20110 21505 20128 21539
rect 20076 21496 20128 21505
rect 22008 21539 22060 21548
rect 22008 21505 22017 21539
rect 22017 21505 22051 21539
rect 22051 21505 22060 21539
rect 22008 21496 22060 21505
rect 23572 21496 23624 21548
rect 24032 21539 24084 21548
rect 24032 21505 24041 21539
rect 24041 21505 24075 21539
rect 24075 21505 24084 21539
rect 24032 21496 24084 21505
rect 24216 21496 24268 21548
rect 25044 21496 25096 21548
rect 26240 21496 26292 21548
rect 27344 21539 27396 21548
rect 27344 21505 27353 21539
rect 27353 21505 27387 21539
rect 27387 21505 27396 21539
rect 27344 21496 27396 21505
rect 28816 21496 28868 21548
rect 31760 21632 31812 21684
rect 32588 21632 32640 21684
rect 35716 21632 35768 21684
rect 30288 21564 30340 21616
rect 29920 21496 29972 21548
rect 31392 21564 31444 21616
rect 33508 21607 33560 21616
rect 32588 21539 32640 21548
rect 27528 21428 27580 21480
rect 28172 21471 28224 21480
rect 28172 21437 28181 21471
rect 28181 21437 28215 21471
rect 28215 21437 28224 21471
rect 28172 21428 28224 21437
rect 28080 21360 28132 21412
rect 28448 21471 28500 21480
rect 28448 21437 28457 21471
rect 28457 21437 28491 21471
rect 28491 21437 28500 21471
rect 28448 21428 28500 21437
rect 28632 21428 28684 21480
rect 28908 21360 28960 21412
rect 23480 21292 23532 21344
rect 25228 21292 25280 21344
rect 25504 21292 25556 21344
rect 26700 21292 26752 21344
rect 30932 21292 30984 21344
rect 32588 21505 32597 21539
rect 32597 21505 32631 21539
rect 32631 21505 32640 21539
rect 32588 21496 32640 21505
rect 33508 21573 33517 21607
rect 33517 21573 33551 21607
rect 33551 21573 33560 21607
rect 33508 21564 33560 21573
rect 34704 21564 34756 21616
rect 35624 21564 35676 21616
rect 36176 21632 36228 21684
rect 37648 21564 37700 21616
rect 32680 21360 32732 21412
rect 34152 21428 34204 21480
rect 36636 21496 36688 21548
rect 34796 21428 34848 21480
rect 35532 21292 35584 21344
rect 35624 21292 35676 21344
rect 36176 21292 36228 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 23572 21088 23624 21140
rect 28172 21088 28224 21140
rect 28356 21020 28408 21072
rect 28632 21020 28684 21072
rect 24308 20952 24360 21004
rect 29736 20952 29788 21004
rect 30012 20952 30064 21004
rect 1768 20927 1820 20936
rect 1768 20893 1777 20927
rect 1777 20893 1811 20927
rect 1811 20893 1820 20927
rect 1768 20884 1820 20893
rect 22008 20884 22060 20936
rect 23572 20884 23624 20936
rect 27712 20884 27764 20936
rect 28632 20927 28684 20936
rect 28632 20893 28641 20927
rect 28641 20893 28675 20927
rect 28675 20893 28684 20927
rect 28632 20884 28684 20893
rect 30564 20927 30616 20936
rect 30564 20893 30598 20927
rect 30598 20893 30616 20927
rect 30564 20884 30616 20893
rect 32404 20884 32456 20936
rect 35532 20884 35584 20936
rect 23480 20816 23532 20868
rect 24860 20859 24912 20868
rect 24860 20825 24894 20859
rect 24894 20825 24912 20859
rect 26700 20859 26752 20868
rect 24860 20816 24912 20825
rect 26700 20825 26734 20859
rect 26734 20825 26752 20859
rect 26700 20816 26752 20825
rect 27528 20816 27580 20868
rect 33140 20816 33192 20868
rect 35992 20816 36044 20868
rect 25136 20748 25188 20800
rect 27988 20748 28040 20800
rect 28540 20791 28592 20800
rect 28540 20757 28549 20791
rect 28549 20757 28583 20791
rect 28583 20757 28592 20791
rect 31668 20791 31720 20800
rect 28540 20748 28592 20757
rect 31668 20757 31677 20791
rect 31677 20757 31711 20791
rect 31711 20757 31720 20791
rect 31668 20748 31720 20757
rect 32496 20748 32548 20800
rect 35256 20748 35308 20800
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 24860 20544 24912 20596
rect 20628 20408 20680 20460
rect 24032 20476 24084 20528
rect 24216 20408 24268 20460
rect 24860 20408 24912 20460
rect 27712 20476 27764 20528
rect 25504 20451 25556 20460
rect 25504 20417 25538 20451
rect 25538 20417 25556 20451
rect 25504 20408 25556 20417
rect 25136 20340 25188 20392
rect 24032 20272 24084 20324
rect 27528 20408 27580 20460
rect 27988 20451 28040 20460
rect 27988 20417 27997 20451
rect 27997 20417 28031 20451
rect 28031 20417 28040 20451
rect 29092 20544 29144 20596
rect 31116 20544 31168 20596
rect 32588 20544 32640 20596
rect 33140 20544 33192 20596
rect 35992 20587 36044 20596
rect 35992 20553 36001 20587
rect 36001 20553 36035 20587
rect 36035 20553 36044 20587
rect 35992 20544 36044 20553
rect 36636 20587 36688 20596
rect 36636 20553 36645 20587
rect 36645 20553 36679 20587
rect 36679 20553 36688 20587
rect 36636 20544 36688 20553
rect 29000 20519 29052 20528
rect 29000 20485 29034 20519
rect 29034 20485 29052 20519
rect 29000 20476 29052 20485
rect 32496 20476 32548 20528
rect 34796 20476 34848 20528
rect 27988 20408 28040 20417
rect 27712 20340 27764 20392
rect 30564 20340 30616 20392
rect 30932 20340 30984 20392
rect 31668 20340 31720 20392
rect 33508 20408 33560 20460
rect 35256 20451 35308 20460
rect 35256 20417 35265 20451
rect 35265 20417 35299 20451
rect 35299 20417 35308 20451
rect 35256 20408 35308 20417
rect 36176 20451 36228 20460
rect 36176 20417 36185 20451
rect 36185 20417 36219 20451
rect 36219 20417 36228 20451
rect 36176 20408 36228 20417
rect 33232 20383 33284 20392
rect 28632 20272 28684 20324
rect 33232 20349 33241 20383
rect 33241 20349 33275 20383
rect 33275 20349 33284 20383
rect 33232 20340 33284 20349
rect 33324 20272 33376 20324
rect 20076 20204 20128 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 28448 20204 28500 20256
rect 28540 20204 28592 20256
rect 31392 20204 31444 20256
rect 33140 20204 33192 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 26240 20043 26292 20052
rect 26240 20009 26249 20043
rect 26249 20009 26283 20043
rect 26283 20009 26292 20043
rect 26240 20000 26292 20009
rect 28356 20043 28408 20052
rect 28356 20009 28365 20043
rect 28365 20009 28399 20043
rect 28399 20009 28408 20043
rect 28356 20000 28408 20009
rect 28632 20043 28684 20052
rect 28632 20009 28641 20043
rect 28641 20009 28675 20043
rect 28675 20009 28684 20043
rect 28632 20000 28684 20009
rect 33232 20000 33284 20052
rect 25780 19932 25832 19984
rect 25596 19864 25648 19916
rect 27988 19864 28040 19916
rect 31668 19864 31720 19916
rect 33508 19864 33560 19916
rect 19432 19796 19484 19848
rect 22192 19839 22244 19848
rect 22192 19805 22201 19839
rect 22201 19805 22235 19839
rect 22235 19805 22244 19839
rect 22192 19796 22244 19805
rect 23848 19839 23900 19848
rect 20352 19728 20404 19780
rect 21640 19728 21692 19780
rect 23848 19805 23857 19839
rect 23857 19805 23891 19839
rect 23891 19805 23900 19839
rect 23848 19796 23900 19805
rect 24032 19839 24084 19848
rect 24032 19805 24041 19839
rect 24041 19805 24075 19839
rect 24075 19805 24084 19839
rect 24032 19796 24084 19805
rect 25136 19839 25188 19848
rect 25136 19805 25145 19839
rect 25145 19805 25179 19839
rect 25179 19805 25188 19839
rect 25136 19796 25188 19805
rect 27344 19796 27396 19848
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 28540 19796 28592 19848
rect 29920 19839 29972 19848
rect 29920 19805 29929 19839
rect 29929 19805 29963 19839
rect 29963 19805 29972 19839
rect 29920 19796 29972 19805
rect 30564 19796 30616 19848
rect 31576 19796 31628 19848
rect 32404 19796 32456 19848
rect 35992 19839 36044 19848
rect 25228 19728 25280 19780
rect 27160 19728 27212 19780
rect 33416 19728 33468 19780
rect 35992 19805 36001 19839
rect 36001 19805 36035 19839
rect 36035 19805 36044 19839
rect 35992 19796 36044 19805
rect 36544 19728 36596 19780
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 22284 19703 22336 19712
rect 22284 19669 22293 19703
rect 22293 19669 22327 19703
rect 22327 19669 22336 19703
rect 22284 19660 22336 19669
rect 23480 19660 23532 19712
rect 25964 19660 26016 19712
rect 29460 19660 29512 19712
rect 30932 19660 30984 19712
rect 34704 19660 34756 19712
rect 35808 19703 35860 19712
rect 35808 19669 35817 19703
rect 35817 19669 35851 19703
rect 35851 19669 35860 19703
rect 35808 19660 35860 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 20352 19499 20404 19508
rect 20352 19465 20361 19499
rect 20361 19465 20395 19499
rect 20395 19465 20404 19499
rect 20352 19456 20404 19465
rect 25596 19499 25648 19508
rect 25596 19465 25605 19499
rect 25605 19465 25639 19499
rect 25639 19465 25648 19499
rect 25596 19456 25648 19465
rect 19432 19388 19484 19440
rect 22284 19431 22336 19440
rect 22284 19397 22318 19431
rect 22318 19397 22336 19431
rect 22284 19388 22336 19397
rect 28264 19456 28316 19508
rect 30472 19456 30524 19508
rect 32680 19456 32732 19508
rect 32864 19456 32916 19508
rect 33600 19499 33652 19508
rect 33600 19465 33609 19499
rect 33609 19465 33643 19499
rect 33643 19465 33652 19499
rect 33600 19456 33652 19465
rect 37004 19456 37056 19508
rect 33140 19388 33192 19440
rect 33232 19431 33284 19440
rect 33232 19397 33241 19431
rect 33241 19397 33275 19431
rect 33275 19397 33284 19431
rect 35808 19431 35860 19440
rect 33232 19388 33284 19397
rect 35808 19397 35842 19431
rect 35842 19397 35860 19431
rect 35808 19388 35860 19397
rect 20536 19363 20588 19372
rect 20168 19252 20220 19304
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 22008 19363 22060 19372
rect 22008 19329 22017 19363
rect 22017 19329 22051 19363
rect 22051 19329 22060 19363
rect 22008 19320 22060 19329
rect 26240 19363 26292 19372
rect 26240 19329 26249 19363
rect 26249 19329 26283 19363
rect 26283 19329 26292 19363
rect 26240 19320 26292 19329
rect 27344 19363 27396 19372
rect 27344 19329 27353 19363
rect 27353 19329 27387 19363
rect 27387 19329 27396 19363
rect 27344 19320 27396 19329
rect 28172 19363 28224 19372
rect 28172 19329 28181 19363
rect 28181 19329 28215 19363
rect 28215 19329 28224 19363
rect 28172 19320 28224 19329
rect 28264 19320 28316 19372
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 29644 19320 29696 19372
rect 30932 19363 30984 19372
rect 30932 19329 30941 19363
rect 30941 19329 30975 19363
rect 30975 19329 30984 19363
rect 30932 19320 30984 19329
rect 31576 19363 31628 19372
rect 31576 19329 31585 19363
rect 31585 19329 31619 19363
rect 31619 19329 31628 19363
rect 31576 19320 31628 19329
rect 32312 19363 32364 19372
rect 32312 19329 32321 19363
rect 32321 19329 32355 19363
rect 32355 19329 32364 19363
rect 32312 19320 32364 19329
rect 32588 19363 32640 19372
rect 32588 19329 32597 19363
rect 32597 19329 32631 19363
rect 32631 19329 32640 19363
rect 32588 19320 32640 19329
rect 34704 19363 34756 19372
rect 34704 19329 34713 19363
rect 34713 19329 34747 19363
rect 34747 19329 34756 19363
rect 34704 19320 34756 19329
rect 37648 19363 37700 19372
rect 37648 19329 37657 19363
rect 37657 19329 37691 19363
rect 37691 19329 37700 19363
rect 37648 19320 37700 19329
rect 20720 19252 20772 19304
rect 21272 19252 21324 19304
rect 24216 19295 24268 19304
rect 24216 19261 24225 19295
rect 24225 19261 24259 19295
rect 24259 19261 24268 19295
rect 24216 19252 24268 19261
rect 28356 19295 28408 19304
rect 28356 19261 28365 19295
rect 28365 19261 28399 19295
rect 28399 19261 28408 19295
rect 28356 19252 28408 19261
rect 31392 19295 31444 19304
rect 31392 19261 31401 19295
rect 31401 19261 31435 19295
rect 31435 19261 31444 19295
rect 31392 19252 31444 19261
rect 33232 19252 33284 19304
rect 35532 19295 35584 19304
rect 35532 19261 35541 19295
rect 35541 19261 35575 19295
rect 35575 19261 35584 19295
rect 35532 19252 35584 19261
rect 19708 19159 19760 19168
rect 19708 19125 19717 19159
rect 19717 19125 19751 19159
rect 19751 19125 19760 19159
rect 19708 19116 19760 19125
rect 20812 19116 20864 19168
rect 21640 19116 21692 19168
rect 22376 19116 22428 19168
rect 27252 19116 27304 19168
rect 28724 19116 28776 19168
rect 29828 19116 29880 19168
rect 29920 19159 29972 19168
rect 29920 19125 29929 19159
rect 29929 19125 29963 19159
rect 29963 19125 29972 19159
rect 32496 19159 32548 19168
rect 29920 19116 29972 19125
rect 32496 19125 32505 19159
rect 32505 19125 32539 19159
rect 32539 19125 32548 19159
rect 32496 19116 32548 19125
rect 33324 19116 33376 19168
rect 34704 19116 34756 19168
rect 36636 19116 36688 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 25964 18955 26016 18964
rect 25964 18921 25973 18955
rect 25973 18921 26007 18955
rect 26007 18921 26016 18955
rect 25964 18912 26016 18921
rect 28816 18955 28868 18964
rect 28816 18921 28825 18955
rect 28825 18921 28859 18955
rect 28859 18921 28868 18955
rect 28816 18912 28868 18921
rect 33416 18955 33468 18964
rect 33416 18921 33425 18955
rect 33425 18921 33459 18955
rect 33459 18921 33468 18955
rect 33416 18912 33468 18921
rect 32404 18776 32456 18828
rect 19432 18708 19484 18760
rect 19708 18708 19760 18760
rect 21272 18708 21324 18760
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 22008 18708 22060 18760
rect 23572 18708 23624 18760
rect 24216 18708 24268 18760
rect 24676 18708 24728 18760
rect 27528 18708 27580 18760
rect 28264 18751 28316 18760
rect 28264 18717 28273 18751
rect 28273 18717 28307 18751
rect 28307 18717 28316 18751
rect 28264 18708 28316 18717
rect 28356 18708 28408 18760
rect 31208 18751 31260 18760
rect 31208 18717 31217 18751
rect 31217 18717 31251 18751
rect 31251 18717 31260 18751
rect 31208 18708 31260 18717
rect 33140 18708 33192 18760
rect 34244 18751 34296 18760
rect 34244 18717 34253 18751
rect 34253 18717 34287 18751
rect 34287 18717 34296 18751
rect 34244 18708 34296 18717
rect 34520 18708 34572 18760
rect 35532 18708 35584 18760
rect 37004 18751 37056 18760
rect 37004 18717 37038 18751
rect 37038 18717 37056 18751
rect 37004 18708 37056 18717
rect 19984 18640 20036 18692
rect 20628 18640 20680 18692
rect 23480 18640 23532 18692
rect 25596 18640 25648 18692
rect 28080 18640 28132 18692
rect 28724 18640 28776 18692
rect 34704 18640 34756 18692
rect 21180 18572 21232 18624
rect 23112 18572 23164 18624
rect 25044 18572 25096 18624
rect 27712 18572 27764 18624
rect 28172 18572 28224 18624
rect 34060 18615 34112 18624
rect 34060 18581 34069 18615
rect 34069 18581 34103 18615
rect 34103 18581 34112 18615
rect 34060 18572 34112 18581
rect 36268 18615 36320 18624
rect 36268 18581 36277 18615
rect 36277 18581 36311 18615
rect 36311 18581 36320 18615
rect 36268 18572 36320 18581
rect 37464 18572 37516 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 20168 18411 20220 18420
rect 20168 18377 20177 18411
rect 20177 18377 20211 18411
rect 20211 18377 20220 18411
rect 20168 18368 20220 18377
rect 20812 18411 20864 18420
rect 20812 18377 20837 18411
rect 20837 18377 20864 18411
rect 20812 18368 20864 18377
rect 22192 18368 22244 18420
rect 23572 18368 23624 18420
rect 25596 18411 25648 18420
rect 25596 18377 25605 18411
rect 25605 18377 25639 18411
rect 25639 18377 25648 18411
rect 25596 18368 25648 18377
rect 28356 18368 28408 18420
rect 28816 18368 28868 18420
rect 33232 18368 33284 18420
rect 35992 18411 36044 18420
rect 35992 18377 36001 18411
rect 36001 18377 36035 18411
rect 36035 18377 36044 18411
rect 35992 18368 36044 18377
rect 21180 18300 21232 18352
rect 19984 18275 20036 18284
rect 19984 18241 19993 18275
rect 19993 18241 20027 18275
rect 20027 18241 20036 18275
rect 22376 18275 22428 18284
rect 19984 18232 20036 18241
rect 22376 18241 22385 18275
rect 22385 18241 22419 18275
rect 22419 18241 22428 18275
rect 22376 18232 22428 18241
rect 22100 18164 22152 18216
rect 24124 18300 24176 18352
rect 23388 18275 23440 18284
rect 23388 18241 23397 18275
rect 23397 18241 23431 18275
rect 23431 18241 23440 18275
rect 23388 18232 23440 18241
rect 25780 18275 25832 18284
rect 25780 18241 25789 18275
rect 25789 18241 25823 18275
rect 25823 18241 25832 18275
rect 25780 18232 25832 18241
rect 25964 18232 26016 18284
rect 27528 18300 27580 18352
rect 34060 18300 34112 18352
rect 34704 18343 34756 18352
rect 34704 18309 34713 18343
rect 34713 18309 34747 18343
rect 34747 18309 34756 18343
rect 34704 18300 34756 18309
rect 27252 18232 27304 18284
rect 29736 18275 29788 18284
rect 29736 18241 29745 18275
rect 29745 18241 29779 18275
rect 29779 18241 29788 18275
rect 29736 18232 29788 18241
rect 29828 18232 29880 18284
rect 32404 18275 32456 18284
rect 32404 18241 32413 18275
rect 32413 18241 32447 18275
rect 32447 18241 32456 18275
rect 32404 18232 32456 18241
rect 20720 18096 20772 18148
rect 21272 18028 21324 18080
rect 24032 18028 24084 18080
rect 25136 18028 25188 18080
rect 25872 18028 25924 18080
rect 31208 18096 31260 18148
rect 34704 18164 34756 18216
rect 35348 18164 35400 18216
rect 36268 18300 36320 18352
rect 35900 18232 35952 18284
rect 37556 18300 37608 18352
rect 37464 18164 37516 18216
rect 34428 18071 34480 18080
rect 34428 18037 34437 18071
rect 34437 18037 34471 18071
rect 34471 18037 34480 18071
rect 34428 18028 34480 18037
rect 36544 18071 36596 18080
rect 36544 18037 36553 18071
rect 36553 18037 36587 18071
rect 36587 18037 36596 18071
rect 36544 18028 36596 18037
rect 36820 18071 36872 18080
rect 36820 18037 36829 18071
rect 36829 18037 36863 18071
rect 36863 18037 36872 18071
rect 36820 18028 36872 18037
rect 36912 18028 36964 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 20720 17824 20772 17876
rect 21640 17756 21692 17808
rect 20444 17663 20496 17672
rect 20444 17629 20453 17663
rect 20453 17629 20487 17663
rect 20487 17629 20496 17663
rect 20444 17620 20496 17629
rect 20720 17620 20772 17672
rect 22652 17620 22704 17672
rect 24032 17824 24084 17876
rect 25964 17867 26016 17876
rect 25964 17833 25973 17867
rect 25973 17833 26007 17867
rect 26007 17833 26016 17867
rect 25964 17824 26016 17833
rect 27344 17824 27396 17876
rect 28080 17824 28132 17876
rect 29828 17824 29880 17876
rect 34244 17824 34296 17876
rect 35348 17824 35400 17876
rect 37648 17824 37700 17876
rect 23112 17663 23164 17672
rect 23112 17629 23121 17663
rect 23121 17629 23155 17663
rect 23155 17629 23164 17663
rect 23112 17620 23164 17629
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 24584 17620 24636 17672
rect 25504 17756 25556 17808
rect 28264 17756 28316 17808
rect 36820 17756 36872 17808
rect 25136 17663 25188 17672
rect 25136 17629 25150 17663
rect 25150 17629 25184 17663
rect 25184 17629 25188 17663
rect 25136 17620 25188 17629
rect 20904 17595 20956 17604
rect 20904 17561 20913 17595
rect 20913 17561 20947 17595
rect 20947 17561 20956 17595
rect 20904 17552 20956 17561
rect 22192 17552 22244 17604
rect 22376 17552 22428 17604
rect 25228 17552 25280 17604
rect 25412 17552 25464 17604
rect 25872 17552 25924 17604
rect 26516 17552 26568 17604
rect 26792 17663 26844 17672
rect 26792 17629 26801 17663
rect 26801 17629 26835 17663
rect 26835 17629 26844 17663
rect 26792 17620 26844 17629
rect 28816 17663 28868 17672
rect 28816 17629 28825 17663
rect 28825 17629 28859 17663
rect 28859 17629 28868 17663
rect 28816 17620 28868 17629
rect 32496 17688 32548 17740
rect 30564 17663 30616 17672
rect 27712 17552 27764 17604
rect 30564 17629 30573 17663
rect 30573 17629 30607 17663
rect 30607 17629 30616 17663
rect 30564 17620 30616 17629
rect 31208 17663 31260 17672
rect 31208 17629 31217 17663
rect 31217 17629 31251 17663
rect 31251 17629 31260 17663
rect 31208 17620 31260 17629
rect 32312 17620 32364 17672
rect 33416 17663 33468 17672
rect 33416 17629 33425 17663
rect 33425 17629 33459 17663
rect 33459 17629 33468 17663
rect 33416 17620 33468 17629
rect 31576 17552 31628 17604
rect 35532 17620 35584 17672
rect 36636 17663 36688 17672
rect 34796 17552 34848 17604
rect 36636 17629 36645 17663
rect 36645 17629 36679 17663
rect 36679 17629 36688 17663
rect 36636 17620 36688 17629
rect 37464 17663 37516 17672
rect 35900 17552 35952 17604
rect 37464 17629 37473 17663
rect 37473 17629 37507 17663
rect 37507 17629 37516 17663
rect 37464 17620 37516 17629
rect 19984 17527 20036 17536
rect 19984 17493 19993 17527
rect 19993 17493 20027 17527
rect 20027 17493 20036 17527
rect 19984 17484 20036 17493
rect 20444 17484 20496 17536
rect 23664 17484 23716 17536
rect 26148 17527 26200 17536
rect 26148 17493 26157 17527
rect 26157 17493 26191 17527
rect 26191 17493 26200 17527
rect 26148 17484 26200 17493
rect 29000 17484 29052 17536
rect 30748 17527 30800 17536
rect 30748 17493 30757 17527
rect 30757 17493 30791 17527
rect 30791 17493 30800 17527
rect 30748 17484 30800 17493
rect 37648 17484 37700 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 23848 17280 23900 17332
rect 24676 17323 24728 17332
rect 24676 17289 24685 17323
rect 24685 17289 24719 17323
rect 24719 17289 24728 17323
rect 24676 17280 24728 17289
rect 25136 17280 25188 17332
rect 25964 17280 26016 17332
rect 28264 17280 28316 17332
rect 19984 17212 20036 17264
rect 23388 17255 23440 17264
rect 23388 17221 23397 17255
rect 23397 17221 23431 17255
rect 23431 17221 23440 17255
rect 23388 17212 23440 17221
rect 25320 17212 25372 17264
rect 27160 17255 27212 17264
rect 27160 17221 27169 17255
rect 27169 17221 27203 17255
rect 27203 17221 27212 17255
rect 27160 17212 27212 17221
rect 27528 17212 27580 17264
rect 19432 17144 19484 17196
rect 22652 17187 22704 17196
rect 22652 17153 22661 17187
rect 22661 17153 22695 17187
rect 22695 17153 22704 17187
rect 22652 17144 22704 17153
rect 23296 17144 23348 17196
rect 26148 17144 26200 17196
rect 26516 17144 26568 17196
rect 27252 17144 27304 17196
rect 28724 17212 28776 17264
rect 30472 17255 30524 17264
rect 30472 17221 30506 17255
rect 30506 17221 30524 17255
rect 30472 17212 30524 17221
rect 32220 17212 32272 17264
rect 32588 17280 32640 17332
rect 32864 17323 32916 17332
rect 32864 17289 32873 17323
rect 32873 17289 32907 17323
rect 32907 17289 32916 17323
rect 32864 17280 32916 17289
rect 34796 17323 34848 17332
rect 34796 17289 34805 17323
rect 34805 17289 34839 17323
rect 34839 17289 34848 17323
rect 34796 17280 34848 17289
rect 35532 17280 35584 17332
rect 32496 17255 32548 17264
rect 32496 17221 32505 17255
rect 32505 17221 32539 17255
rect 32539 17221 32548 17255
rect 32496 17212 32548 17221
rect 28448 17144 28500 17196
rect 29736 17144 29788 17196
rect 30196 17187 30248 17196
rect 30196 17153 30205 17187
rect 30205 17153 30239 17187
rect 30239 17153 30248 17187
rect 30196 17144 30248 17153
rect 33232 17212 33284 17264
rect 34428 17212 34480 17264
rect 37280 17212 37332 17264
rect 35440 17187 35492 17196
rect 24952 17076 25004 17128
rect 24860 17008 24912 17060
rect 32312 17076 32364 17128
rect 35440 17153 35449 17187
rect 35449 17153 35483 17187
rect 35483 17153 35492 17187
rect 35440 17144 35492 17153
rect 37648 17187 37700 17196
rect 32496 17008 32548 17060
rect 20168 16940 20220 16992
rect 20444 16940 20496 16992
rect 20628 16940 20680 16992
rect 25596 16983 25648 16992
rect 25596 16949 25605 16983
rect 25605 16949 25639 16983
rect 25639 16949 25648 16983
rect 25596 16940 25648 16949
rect 27344 16940 27396 16992
rect 36268 17076 36320 17128
rect 36360 17008 36412 17060
rect 37648 17153 37657 17187
rect 37657 17153 37691 17187
rect 37691 17153 37700 17187
rect 37648 17144 37700 17153
rect 34520 16940 34572 16992
rect 35348 16940 35400 16992
rect 36544 16983 36596 16992
rect 36544 16949 36553 16983
rect 36553 16949 36587 16983
rect 36587 16949 36596 16983
rect 36544 16940 36596 16949
rect 37188 16940 37240 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 22192 16736 22244 16788
rect 20444 16668 20496 16720
rect 20628 16668 20680 16720
rect 21272 16668 21324 16720
rect 20260 16575 20312 16584
rect 20260 16541 20269 16575
rect 20269 16541 20303 16575
rect 20303 16541 20312 16575
rect 20260 16532 20312 16541
rect 20720 16532 20772 16584
rect 22192 16575 22244 16584
rect 21180 16464 21232 16516
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 22192 16541 22201 16575
rect 22201 16541 22235 16575
rect 22235 16541 22244 16575
rect 22192 16532 22244 16541
rect 23480 16668 23532 16720
rect 24584 16736 24636 16788
rect 28448 16736 28500 16788
rect 30196 16736 30248 16788
rect 33416 16779 33468 16788
rect 22836 16532 22888 16584
rect 23664 16600 23716 16652
rect 24676 16600 24728 16652
rect 30196 16643 30248 16652
rect 30196 16609 30205 16643
rect 30205 16609 30239 16643
rect 30239 16609 30248 16643
rect 30196 16600 30248 16609
rect 33416 16745 33425 16779
rect 33425 16745 33459 16779
rect 33459 16745 33468 16779
rect 33416 16736 33468 16745
rect 34520 16736 34572 16788
rect 33968 16668 34020 16720
rect 36268 16711 36320 16720
rect 36268 16677 36277 16711
rect 36277 16677 36311 16711
rect 36311 16677 36320 16711
rect 36268 16668 36320 16677
rect 36912 16643 36964 16652
rect 36912 16609 36921 16643
rect 36921 16609 36955 16643
rect 36955 16609 36964 16643
rect 36912 16600 36964 16609
rect 24952 16575 25004 16584
rect 24952 16541 24961 16575
rect 24961 16541 24995 16575
rect 24995 16541 25004 16575
rect 24952 16532 25004 16541
rect 25136 16575 25188 16584
rect 25136 16541 25145 16575
rect 25145 16541 25179 16575
rect 25179 16541 25188 16575
rect 25136 16532 25188 16541
rect 22744 16439 22796 16448
rect 22744 16405 22753 16439
rect 22753 16405 22787 16439
rect 22787 16405 22796 16439
rect 22744 16396 22796 16405
rect 23112 16464 23164 16516
rect 23480 16507 23532 16516
rect 23480 16473 23489 16507
rect 23489 16473 23523 16507
rect 23523 16473 23532 16507
rect 25320 16575 25372 16584
rect 25320 16541 25329 16575
rect 25329 16541 25363 16575
rect 25363 16541 25372 16575
rect 25320 16532 25372 16541
rect 25504 16575 25556 16584
rect 25504 16541 25513 16575
rect 25513 16541 25547 16575
rect 25547 16541 25556 16575
rect 25504 16532 25556 16541
rect 28908 16532 28960 16584
rect 23480 16464 23532 16473
rect 25412 16464 25464 16516
rect 27160 16464 27212 16516
rect 34796 16532 34848 16584
rect 37188 16575 37240 16584
rect 37188 16541 37222 16575
rect 37222 16541 37240 16575
rect 37188 16532 37240 16541
rect 27528 16396 27580 16448
rect 30564 16464 30616 16516
rect 30840 16464 30892 16516
rect 35348 16464 35400 16516
rect 29092 16439 29144 16448
rect 29092 16405 29101 16439
rect 29101 16405 29135 16439
rect 29135 16405 29144 16439
rect 29092 16396 29144 16405
rect 32128 16396 32180 16448
rect 34336 16439 34388 16448
rect 34336 16405 34345 16439
rect 34345 16405 34379 16439
rect 34379 16405 34388 16439
rect 34336 16396 34388 16405
rect 37188 16396 37240 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 20628 16192 20680 16244
rect 20168 16124 20220 16176
rect 20076 16056 20128 16108
rect 22744 16192 22796 16244
rect 24952 16192 25004 16244
rect 27160 16235 27212 16244
rect 27160 16201 27169 16235
rect 27169 16201 27203 16235
rect 27203 16201 27212 16235
rect 27160 16192 27212 16201
rect 30564 16235 30616 16244
rect 30564 16201 30573 16235
rect 30573 16201 30607 16235
rect 30607 16201 30616 16235
rect 30564 16192 30616 16201
rect 21272 16124 21324 16176
rect 25596 16124 25648 16176
rect 20904 16099 20956 16108
rect 20904 16065 20911 16099
rect 20911 16065 20956 16099
rect 20904 16056 20956 16065
rect 20444 15988 20496 16040
rect 21180 16099 21232 16108
rect 21180 16065 21194 16099
rect 21194 16065 21228 16099
rect 21228 16065 21232 16099
rect 21180 16056 21232 16065
rect 22100 16056 22152 16108
rect 22376 16099 22428 16108
rect 22376 16065 22385 16099
rect 22385 16065 22419 16099
rect 22419 16065 22428 16099
rect 22376 16056 22428 16065
rect 23572 16056 23624 16108
rect 25136 16056 25188 16108
rect 25872 16056 25924 16108
rect 29092 16124 29144 16176
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 27528 16056 27580 16108
rect 28724 16099 28776 16108
rect 28724 16065 28733 16099
rect 28733 16065 28767 16099
rect 28767 16065 28776 16099
rect 28724 16056 28776 16065
rect 28816 16056 28868 16108
rect 30748 16099 30800 16108
rect 30748 16065 30757 16099
rect 30757 16065 30791 16099
rect 30791 16065 30800 16099
rect 30748 16056 30800 16065
rect 31576 16099 31628 16108
rect 31576 16065 31585 16099
rect 31585 16065 31619 16099
rect 31619 16065 31628 16099
rect 31576 16056 31628 16065
rect 32864 16099 32916 16108
rect 32864 16065 32873 16099
rect 32873 16065 32907 16099
rect 32907 16065 32916 16099
rect 32864 16056 32916 16065
rect 33232 16192 33284 16244
rect 35440 16192 35492 16244
rect 36268 16192 36320 16244
rect 37556 16192 37608 16244
rect 36544 16167 36596 16176
rect 36544 16133 36553 16167
rect 36553 16133 36587 16167
rect 36587 16133 36596 16167
rect 36544 16124 36596 16133
rect 37188 16124 37240 16176
rect 33324 16056 33376 16108
rect 34336 16056 34388 16108
rect 35900 16056 35952 16108
rect 20996 15920 21048 15972
rect 19340 15852 19392 15904
rect 20260 15852 20312 15904
rect 25320 15920 25372 15972
rect 25412 15920 25464 15972
rect 26240 15852 26292 15904
rect 27896 15852 27948 15904
rect 32128 15988 32180 16040
rect 31484 15920 31536 15972
rect 33968 15988 34020 16040
rect 37280 16056 37332 16108
rect 37648 16099 37700 16108
rect 37648 16065 37657 16099
rect 37657 16065 37691 16099
rect 37691 16065 37700 16099
rect 37648 16056 37700 16065
rect 34796 15920 34848 15972
rect 36176 15920 36228 15972
rect 36360 15963 36412 15972
rect 36360 15929 36369 15963
rect 36369 15929 36403 15963
rect 36403 15929 36412 15963
rect 36360 15920 36412 15929
rect 29368 15852 29420 15904
rect 30932 15852 30984 15904
rect 32680 15895 32732 15904
rect 32680 15861 32689 15895
rect 32689 15861 32723 15895
rect 32723 15861 32732 15895
rect 32680 15852 32732 15861
rect 33140 15895 33192 15904
rect 33140 15861 33149 15895
rect 33149 15861 33183 15895
rect 33183 15861 33192 15895
rect 33140 15852 33192 15861
rect 38292 15852 38344 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1860 15648 1912 15700
rect 20444 15691 20496 15700
rect 20444 15657 20453 15691
rect 20453 15657 20487 15691
rect 20487 15657 20496 15691
rect 20444 15648 20496 15657
rect 20904 15648 20956 15700
rect 22836 15648 22888 15700
rect 23112 15691 23164 15700
rect 23112 15657 23121 15691
rect 23121 15657 23155 15691
rect 23155 15657 23164 15691
rect 23112 15648 23164 15657
rect 23480 15648 23532 15700
rect 27804 15648 27856 15700
rect 28816 15648 28868 15700
rect 29092 15648 29144 15700
rect 30380 15648 30432 15700
rect 30840 15648 30892 15700
rect 33232 15691 33284 15700
rect 33232 15657 33241 15691
rect 33241 15657 33275 15691
rect 33275 15657 33284 15691
rect 33232 15648 33284 15657
rect 36176 15648 36228 15700
rect 22376 15580 22428 15632
rect 21180 15444 21232 15496
rect 22100 15487 22152 15496
rect 22100 15453 22109 15487
rect 22109 15453 22143 15487
rect 22143 15453 22152 15487
rect 22100 15444 22152 15453
rect 22652 15444 22704 15496
rect 23664 15444 23716 15496
rect 25320 15444 25372 15496
rect 27252 15512 27304 15564
rect 27896 15512 27948 15564
rect 21456 15376 21508 15428
rect 25228 15376 25280 15428
rect 25872 15376 25924 15428
rect 27528 15376 27580 15428
rect 27712 15487 27764 15496
rect 27712 15453 27721 15487
rect 27721 15453 27755 15487
rect 27755 15453 27764 15487
rect 27712 15444 27764 15453
rect 28540 15444 28592 15496
rect 29092 15487 29144 15496
rect 29092 15453 29101 15487
rect 29101 15453 29135 15487
rect 29135 15453 29144 15487
rect 29092 15444 29144 15453
rect 35900 15580 35952 15632
rect 30932 15487 30984 15496
rect 30932 15453 30941 15487
rect 30941 15453 30975 15487
rect 30975 15453 30984 15487
rect 30932 15444 30984 15453
rect 31484 15487 31536 15496
rect 31484 15453 31493 15487
rect 31493 15453 31527 15487
rect 31527 15453 31536 15487
rect 31484 15444 31536 15453
rect 33140 15512 33192 15564
rect 33324 15555 33376 15564
rect 33324 15521 33333 15555
rect 33333 15521 33367 15555
rect 33367 15521 33376 15555
rect 33324 15512 33376 15521
rect 34796 15512 34848 15564
rect 33048 15487 33100 15496
rect 33048 15453 33057 15487
rect 33057 15453 33091 15487
rect 33091 15453 33100 15487
rect 33048 15444 33100 15453
rect 36176 15487 36228 15496
rect 36176 15453 36185 15487
rect 36185 15453 36219 15487
rect 36219 15453 36228 15487
rect 36176 15444 36228 15453
rect 36912 15555 36964 15564
rect 36912 15521 36921 15555
rect 36921 15521 36955 15555
rect 36955 15521 36964 15555
rect 36912 15512 36964 15521
rect 37648 15444 37700 15496
rect 21364 15308 21416 15360
rect 27620 15351 27672 15360
rect 27620 15317 27629 15351
rect 27629 15317 27663 15351
rect 27663 15317 27672 15351
rect 27620 15308 27672 15317
rect 28908 15308 28960 15360
rect 29368 15308 29420 15360
rect 30656 15308 30708 15360
rect 38108 15376 38160 15428
rect 34888 15351 34940 15360
rect 34888 15317 34897 15351
rect 34897 15317 34931 15351
rect 34931 15317 34940 15351
rect 34888 15308 34940 15317
rect 37648 15308 37700 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 22100 15104 22152 15156
rect 22744 15104 22796 15156
rect 25320 15147 25372 15156
rect 25320 15113 25329 15147
rect 25329 15113 25363 15147
rect 25363 15113 25372 15147
rect 25320 15104 25372 15113
rect 25504 15104 25556 15156
rect 19432 14968 19484 15020
rect 21272 14968 21324 15020
rect 23572 15036 23624 15088
rect 22928 14968 22980 15020
rect 24676 15036 24728 15088
rect 25872 15079 25924 15088
rect 25872 15045 25881 15079
rect 25881 15045 25915 15079
rect 25915 15045 25924 15079
rect 25872 15036 25924 15045
rect 24032 14968 24084 15020
rect 26332 14968 26384 15020
rect 26424 15011 26476 15020
rect 26424 14977 26433 15011
rect 26433 14977 26467 15011
rect 26467 14977 26476 15011
rect 27712 15104 27764 15156
rect 31392 15104 31444 15156
rect 33140 15147 33192 15156
rect 33140 15113 33149 15147
rect 33149 15113 33183 15147
rect 33183 15113 33192 15147
rect 33140 15104 33192 15113
rect 27528 15079 27580 15088
rect 27528 15045 27537 15079
rect 27537 15045 27571 15079
rect 27571 15045 27580 15079
rect 27528 15036 27580 15045
rect 26424 14968 26476 14977
rect 27620 15011 27672 15020
rect 27620 14977 27629 15011
rect 27629 14977 27663 15011
rect 27663 14977 27672 15011
rect 27620 14968 27672 14977
rect 28908 15011 28960 15020
rect 28908 14977 28917 15011
rect 28917 14977 28951 15011
rect 28951 14977 28960 15011
rect 28908 14968 28960 14977
rect 29368 14968 29420 15020
rect 30012 14968 30064 15020
rect 33048 14968 33100 15020
rect 36636 15104 36688 15156
rect 38108 15147 38160 15156
rect 38108 15113 38117 15147
rect 38117 15113 38151 15147
rect 38151 15113 38160 15147
rect 38108 15104 38160 15113
rect 34888 14968 34940 15020
rect 35900 15036 35952 15088
rect 36912 15036 36964 15088
rect 35532 14968 35584 15020
rect 37648 15011 37700 15020
rect 37648 14977 37657 15011
rect 37657 14977 37691 15011
rect 37691 14977 37700 15011
rect 37648 14968 37700 14977
rect 38292 15011 38344 15020
rect 38292 14977 38301 15011
rect 38301 14977 38335 15011
rect 38335 14977 38344 15011
rect 38292 14968 38344 14977
rect 28724 14900 28776 14952
rect 32588 14900 32640 14952
rect 28080 14832 28132 14884
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 27344 14807 27396 14816
rect 27344 14773 27353 14807
rect 27353 14773 27387 14807
rect 27387 14773 27396 14807
rect 27344 14764 27396 14773
rect 28908 14764 28960 14816
rect 32680 14764 32732 14816
rect 37464 14807 37516 14816
rect 37464 14773 37473 14807
rect 37473 14773 37507 14807
rect 37507 14773 37516 14807
rect 37464 14764 37516 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 21272 14603 21324 14612
rect 21272 14569 21281 14603
rect 21281 14569 21315 14603
rect 21315 14569 21324 14603
rect 21272 14560 21324 14569
rect 24032 14560 24084 14612
rect 27620 14603 27672 14612
rect 27620 14569 27629 14603
rect 27629 14569 27663 14603
rect 27663 14569 27672 14603
rect 27620 14560 27672 14569
rect 27804 14603 27856 14612
rect 27804 14569 27813 14603
rect 27813 14569 27847 14603
rect 27847 14569 27856 14603
rect 27804 14560 27856 14569
rect 30012 14603 30064 14612
rect 30012 14569 30021 14603
rect 30021 14569 30055 14603
rect 30055 14569 30064 14603
rect 30012 14560 30064 14569
rect 32588 14603 32640 14612
rect 32588 14569 32597 14603
rect 32597 14569 32631 14603
rect 32631 14569 32640 14603
rect 32588 14560 32640 14569
rect 32956 14560 33008 14612
rect 35532 14560 35584 14612
rect 37280 14603 37332 14612
rect 37280 14569 37289 14603
rect 37289 14569 37323 14603
rect 37323 14569 37332 14603
rect 37280 14560 37332 14569
rect 19432 14467 19484 14476
rect 19432 14433 19441 14467
rect 19441 14433 19475 14467
rect 19475 14433 19484 14467
rect 19432 14424 19484 14433
rect 21548 14399 21600 14408
rect 21548 14365 21557 14399
rect 21557 14365 21591 14399
rect 21591 14365 21600 14399
rect 21548 14356 21600 14365
rect 20444 14288 20496 14340
rect 20076 14220 20128 14272
rect 21364 14288 21416 14340
rect 20812 14263 20864 14272
rect 20812 14229 20821 14263
rect 20821 14229 20855 14263
rect 20855 14229 20864 14263
rect 20812 14220 20864 14229
rect 21272 14220 21324 14272
rect 23572 14356 23624 14408
rect 24124 14424 24176 14476
rect 24676 14424 24728 14476
rect 28724 14424 28776 14476
rect 23940 14288 23992 14340
rect 25780 14356 25832 14408
rect 27988 14356 28040 14408
rect 30196 14399 30248 14408
rect 25228 14331 25280 14340
rect 25228 14297 25262 14331
rect 25262 14297 25280 14331
rect 25228 14288 25280 14297
rect 27528 14288 27580 14340
rect 27712 14288 27764 14340
rect 27896 14288 27948 14340
rect 30196 14365 30205 14399
rect 30205 14365 30239 14399
rect 30239 14365 30248 14399
rect 30196 14356 30248 14365
rect 30656 14356 30708 14408
rect 33048 14399 33100 14408
rect 33048 14365 33057 14399
rect 33057 14365 33091 14399
rect 33091 14365 33100 14399
rect 33048 14356 33100 14365
rect 35900 14467 35952 14476
rect 35900 14433 35909 14467
rect 35909 14433 35943 14467
rect 35943 14433 35952 14467
rect 35900 14424 35952 14433
rect 35440 14399 35492 14408
rect 35440 14365 35449 14399
rect 35449 14365 35483 14399
rect 35483 14365 35492 14399
rect 35440 14356 35492 14365
rect 37464 14356 37516 14408
rect 28908 14288 28960 14340
rect 26332 14263 26384 14272
rect 26332 14229 26341 14263
rect 26341 14229 26375 14263
rect 26375 14229 26384 14263
rect 26332 14220 26384 14229
rect 29000 14220 29052 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 20444 14059 20496 14068
rect 20444 14025 20453 14059
rect 20453 14025 20487 14059
rect 20487 14025 20496 14059
rect 20444 14016 20496 14025
rect 22928 14059 22980 14068
rect 22928 14025 22937 14059
rect 22937 14025 22971 14059
rect 22971 14025 22980 14059
rect 22928 14016 22980 14025
rect 24124 14016 24176 14068
rect 25228 14016 25280 14068
rect 19524 13880 19576 13932
rect 19892 13923 19944 13932
rect 19892 13889 19901 13923
rect 19901 13889 19935 13923
rect 19935 13889 19944 13923
rect 19892 13880 19944 13889
rect 19432 13812 19484 13864
rect 20076 13923 20128 13932
rect 20076 13889 20085 13923
rect 20085 13889 20119 13923
rect 20119 13889 20128 13923
rect 20076 13880 20128 13889
rect 20444 13880 20496 13932
rect 20720 13880 20772 13932
rect 21364 13948 21416 14000
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 22376 13923 22428 13932
rect 22376 13889 22385 13923
rect 22385 13889 22419 13923
rect 22419 13889 22428 13923
rect 22376 13880 22428 13889
rect 23940 13948 23992 14000
rect 27896 14016 27948 14068
rect 22744 13923 22796 13932
rect 22744 13889 22753 13923
rect 22753 13889 22787 13923
rect 22787 13889 22796 13923
rect 22744 13880 22796 13889
rect 23756 13923 23808 13932
rect 23756 13889 23765 13923
rect 23765 13889 23799 13923
rect 23799 13889 23808 13923
rect 23756 13880 23808 13889
rect 26424 13948 26476 14000
rect 21180 13855 21232 13864
rect 21180 13821 21189 13855
rect 21189 13821 21223 13855
rect 21223 13821 21232 13855
rect 21180 13812 21232 13821
rect 22008 13812 22060 13864
rect 22468 13855 22520 13864
rect 19800 13676 19852 13728
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 24860 13812 24912 13864
rect 25596 13923 25648 13932
rect 25596 13889 25605 13923
rect 25605 13889 25639 13923
rect 25639 13889 25648 13923
rect 25596 13880 25648 13889
rect 25780 13923 25832 13932
rect 25780 13889 25789 13923
rect 25789 13889 25823 13923
rect 25823 13889 25832 13923
rect 28080 13948 28132 14000
rect 35440 14016 35492 14068
rect 25780 13880 25832 13889
rect 26332 13812 26384 13864
rect 28632 13880 28684 13932
rect 28724 13880 28776 13932
rect 29184 13948 29236 14000
rect 29092 13923 29144 13932
rect 29092 13889 29126 13923
rect 29126 13889 29144 13923
rect 29092 13880 29144 13889
rect 38108 13880 38160 13932
rect 35808 13855 35860 13864
rect 35808 13821 35817 13855
rect 35817 13821 35851 13855
rect 35851 13821 35860 13855
rect 35808 13812 35860 13821
rect 23848 13719 23900 13728
rect 23848 13685 23857 13719
rect 23857 13685 23891 13719
rect 23891 13685 23900 13719
rect 23848 13676 23900 13685
rect 28356 13676 28408 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19892 13472 19944 13524
rect 19524 13404 19576 13456
rect 20628 13472 20680 13524
rect 21272 13515 21324 13524
rect 21272 13481 21281 13515
rect 21281 13481 21315 13515
rect 21315 13481 21324 13515
rect 21272 13472 21324 13481
rect 22468 13472 22520 13524
rect 25596 13472 25648 13524
rect 29092 13472 29144 13524
rect 30196 13472 30248 13524
rect 20720 13336 20772 13388
rect 22100 13336 22152 13388
rect 27344 13404 27396 13456
rect 27988 13447 28040 13456
rect 27436 13336 27488 13388
rect 19800 13311 19852 13320
rect 19800 13277 19809 13311
rect 19809 13277 19843 13311
rect 19843 13277 19852 13311
rect 19800 13268 19852 13277
rect 20444 13311 20496 13320
rect 20444 13277 20453 13311
rect 20453 13277 20487 13311
rect 20487 13277 20496 13311
rect 20444 13268 20496 13277
rect 20812 13268 20864 13320
rect 20904 13268 20956 13320
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 22468 13268 22520 13320
rect 22284 13200 22336 13252
rect 23848 13268 23900 13320
rect 23940 13311 23992 13320
rect 23940 13277 23949 13311
rect 23949 13277 23983 13311
rect 23983 13277 23992 13311
rect 23940 13268 23992 13277
rect 25964 13311 26016 13320
rect 24676 13200 24728 13252
rect 25964 13277 25973 13311
rect 25973 13277 26007 13311
rect 26007 13277 26016 13311
rect 25964 13268 26016 13277
rect 26700 13311 26752 13320
rect 26700 13277 26709 13311
rect 26709 13277 26743 13311
rect 26743 13277 26752 13311
rect 26700 13268 26752 13277
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 27988 13413 27997 13447
rect 27997 13413 28031 13447
rect 28031 13413 28040 13447
rect 27988 13404 28040 13413
rect 29000 13404 29052 13456
rect 26792 13268 26844 13277
rect 28632 13268 28684 13320
rect 28908 13311 28960 13320
rect 28908 13277 28917 13311
rect 28917 13277 28951 13311
rect 28951 13277 28960 13311
rect 28908 13268 28960 13277
rect 32772 13336 32824 13388
rect 35808 13336 35860 13388
rect 29184 13311 29236 13320
rect 29184 13277 29193 13311
rect 29193 13277 29227 13311
rect 29227 13277 29236 13311
rect 29184 13268 29236 13277
rect 29644 13268 29696 13320
rect 28264 13200 28316 13252
rect 23664 13132 23716 13184
rect 24860 13132 24912 13184
rect 27252 13132 27304 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 20720 12928 20772 12980
rect 22376 12971 22428 12980
rect 22376 12937 22385 12971
rect 22385 12937 22419 12971
rect 22419 12937 22428 12971
rect 22376 12928 22428 12937
rect 23756 12928 23808 12980
rect 24676 12971 24728 12980
rect 24676 12937 24685 12971
rect 24685 12937 24719 12971
rect 24719 12937 24728 12971
rect 24676 12928 24728 12937
rect 28264 12971 28316 12980
rect 28264 12937 28273 12971
rect 28273 12937 28307 12971
rect 28307 12937 28316 12971
rect 28264 12928 28316 12937
rect 28080 12860 28132 12912
rect 20260 12835 20312 12844
rect 20260 12801 20269 12835
rect 20269 12801 20303 12835
rect 20303 12801 20312 12835
rect 20260 12792 20312 12801
rect 22284 12835 22336 12844
rect 22284 12801 22293 12835
rect 22293 12801 22327 12835
rect 22327 12801 22336 12835
rect 22284 12792 22336 12801
rect 22468 12835 22520 12844
rect 22468 12801 22477 12835
rect 22477 12801 22511 12835
rect 22511 12801 22520 12835
rect 22468 12792 22520 12801
rect 22744 12792 22796 12844
rect 23664 12792 23716 12844
rect 24032 12792 24084 12844
rect 24768 12835 24820 12844
rect 20536 12767 20588 12776
rect 20536 12733 20545 12767
rect 20545 12733 20579 12767
rect 20579 12733 20588 12767
rect 20536 12724 20588 12733
rect 22100 12656 22152 12708
rect 23388 12724 23440 12776
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 26332 12792 26384 12844
rect 27436 12792 27488 12844
rect 28356 12835 28408 12844
rect 28356 12801 28365 12835
rect 28365 12801 28399 12835
rect 28399 12801 28408 12835
rect 28356 12792 28408 12801
rect 23940 12656 23992 12708
rect 27252 12724 27304 12776
rect 26240 12656 26292 12708
rect 26332 12699 26384 12708
rect 26332 12665 26341 12699
rect 26341 12665 26375 12699
rect 26375 12665 26384 12699
rect 26332 12656 26384 12665
rect 20444 12631 20496 12640
rect 20444 12597 20453 12631
rect 20453 12597 20487 12631
rect 20487 12597 20496 12631
rect 20444 12588 20496 12597
rect 23480 12588 23532 12640
rect 26424 12631 26476 12640
rect 26424 12597 26433 12631
rect 26433 12597 26467 12631
rect 26467 12597 26476 12631
rect 26424 12588 26476 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 20260 12384 20312 12436
rect 20536 12384 20588 12436
rect 20904 12359 20956 12368
rect 20904 12325 20913 12359
rect 20913 12325 20947 12359
rect 20947 12325 20956 12359
rect 20904 12316 20956 12325
rect 24768 12384 24820 12436
rect 27344 12427 27396 12436
rect 27344 12393 27353 12427
rect 27353 12393 27387 12427
rect 27387 12393 27396 12427
rect 27344 12384 27396 12393
rect 19432 12180 19484 12232
rect 20444 12248 20496 12300
rect 22468 12316 22520 12368
rect 22100 12291 22152 12300
rect 20812 12180 20864 12232
rect 22100 12257 22109 12291
rect 22109 12257 22143 12291
rect 22143 12257 22152 12291
rect 22100 12248 22152 12257
rect 24032 12316 24084 12368
rect 26240 12316 26292 12368
rect 26516 12316 26568 12368
rect 21456 12180 21508 12232
rect 22744 12180 22796 12232
rect 23296 12180 23348 12232
rect 23480 12223 23532 12232
rect 23480 12189 23489 12223
rect 23489 12189 23523 12223
rect 23523 12189 23532 12223
rect 26792 12248 26844 12300
rect 23480 12180 23532 12189
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 27252 12223 27304 12232
rect 26424 12180 26476 12189
rect 27252 12189 27261 12223
rect 27261 12189 27295 12223
rect 27295 12189 27304 12223
rect 27252 12180 27304 12189
rect 26700 12112 26752 12164
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 20812 11883 20864 11892
rect 20812 11849 20821 11883
rect 20821 11849 20855 11883
rect 20855 11849 20864 11883
rect 20812 11840 20864 11849
rect 24032 11883 24084 11892
rect 24032 11849 24041 11883
rect 24041 11849 24075 11883
rect 24075 11849 24084 11883
rect 24032 11840 24084 11849
rect 20260 11704 20312 11756
rect 23664 11747 23716 11756
rect 23664 11713 23673 11747
rect 23673 11713 23707 11747
rect 23707 11713 23716 11747
rect 23664 11704 23716 11713
rect 23940 11636 23992 11688
rect 20536 11543 20588 11552
rect 20536 11509 20545 11543
rect 20545 11509 20579 11543
rect 20579 11509 20588 11543
rect 20536 11500 20588 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 29920 8916 29972 8968
rect 38200 8823 38252 8832
rect 38200 8789 38209 8823
rect 38209 8789 38243 8823
rect 38243 8789 38252 8823
rect 38200 8780 38252 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 29644 2592 29696 2644
rect 38108 2635 38160 2644
rect 38108 2601 38117 2635
rect 38117 2601 38151 2635
rect 38151 2601 38160 2635
rect 38108 2592 38160 2601
rect 1860 2499 1912 2508
rect 1860 2465 1869 2499
rect 1869 2465 1903 2499
rect 1903 2465 1912 2499
rect 1860 2456 1912 2465
rect 20 2388 72 2440
rect 9680 2388 9732 2440
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 29000 2388 29052 2440
rect 38660 2388 38712 2440
rect 19340 2252 19392 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 662 39200 718 39800
rect 10322 39200 10378 39800
rect 19982 39200 20038 39800
rect 29642 39200 29698 39800
rect 39302 39200 39358 39800
rect 676 37262 704 39200
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 10336 37262 10364 39200
rect 19996 37262 20024 39200
rect 29656 37466 29684 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 39316 37466 39344 39200
rect 29644 37460 29696 37466
rect 29644 37402 29696 37408
rect 39304 37460 39356 37466
rect 39304 37402 39356 37408
rect 664 37256 716 37262
rect 664 37198 716 37204
rect 10324 37256 10376 37262
rect 10324 37198 10376 37204
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 32312 37256 32364 37262
rect 32312 37198 32364 37204
rect 1584 37120 1636 37126
rect 1584 37062 1636 37068
rect 10600 37120 10652 37126
rect 10600 37062 10652 37068
rect 24492 37120 24544 37126
rect 24492 37062 24544 37068
rect 1596 31822 1624 37062
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 1584 31816 1636 31822
rect 1584 31758 1636 31764
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 1584 30728 1636 30734
rect 1584 30670 1636 30676
rect 1766 30696 1822 30705
rect 1596 29578 1624 30670
rect 1766 30631 1822 30640
rect 1780 30598 1808 30631
rect 1768 30592 1820 30598
rect 1768 30534 1820 30540
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 1584 29572 1636 29578
rect 1584 29514 1636 29520
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 10612 28218 10640 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23492 33046 23520 33322
rect 23480 33040 23532 33046
rect 23480 32982 23532 32988
rect 23756 33040 23808 33046
rect 23756 32982 23808 32988
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 23768 32366 23796 32982
rect 23860 32910 23888 33798
rect 24032 33516 24084 33522
rect 24032 33458 24084 33464
rect 23940 33448 23992 33454
rect 23940 33390 23992 33396
rect 23952 32910 23980 33390
rect 23848 32904 23900 32910
rect 23848 32846 23900 32852
rect 23940 32904 23992 32910
rect 23940 32846 23992 32852
rect 24044 32774 24072 33458
rect 24032 32768 24084 32774
rect 24032 32710 24084 32716
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 21272 32224 21324 32230
rect 21272 32166 21324 32172
rect 21284 31890 21312 32166
rect 24044 31958 24072 32710
rect 24216 32292 24268 32298
rect 24216 32234 24268 32240
rect 24032 31952 24084 31958
rect 24032 31894 24084 31900
rect 21272 31884 21324 31890
rect 21272 31826 21324 31832
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 20076 31340 20128 31346
rect 20076 31282 20128 31288
rect 19432 31272 19484 31278
rect 19432 31214 19484 31220
rect 17408 30932 17460 30938
rect 17408 30874 17460 30880
rect 17040 30728 17092 30734
rect 17040 30670 17092 30676
rect 16580 30184 16632 30190
rect 16580 30126 16632 30132
rect 16488 29640 16540 29646
rect 16592 29628 16620 30126
rect 17052 29850 17080 30670
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17132 30252 17184 30258
rect 17132 30194 17184 30200
rect 17040 29844 17092 29850
rect 17040 29786 17092 29792
rect 16540 29600 16620 29628
rect 16488 29582 16540 29588
rect 10600 28212 10652 28218
rect 10600 28154 10652 28160
rect 16592 27878 16620 29600
rect 17052 29170 17080 29786
rect 17144 29714 17172 30194
rect 17132 29708 17184 29714
rect 17132 29650 17184 29656
rect 17236 29646 17264 30534
rect 17420 30054 17448 30874
rect 18604 30728 18656 30734
rect 18604 30670 18656 30676
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 17408 30048 17460 30054
rect 17408 29990 17460 29996
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 17316 29708 17368 29714
rect 17316 29650 17368 29656
rect 17224 29640 17276 29646
rect 17224 29582 17276 29588
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17328 29034 17356 29650
rect 17420 29170 17448 29990
rect 18064 29782 18092 29990
rect 18052 29776 18104 29782
rect 18052 29718 18104 29724
rect 18524 29238 18552 30194
rect 18616 29646 18644 30670
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19352 30326 19380 30534
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19444 30258 19472 31214
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19616 30388 19668 30394
rect 19616 30330 19668 30336
rect 19524 30320 19576 30326
rect 19524 30262 19576 30268
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 18880 30184 18932 30190
rect 18880 30126 18932 30132
rect 19064 30184 19116 30190
rect 19116 30144 19380 30172
rect 19064 30126 19116 30132
rect 18892 29850 18920 30126
rect 18880 29844 18932 29850
rect 18880 29786 18932 29792
rect 18800 29714 19104 29730
rect 18788 29708 19104 29714
rect 18840 29702 19104 29708
rect 18788 29650 18840 29656
rect 19076 29646 19104 29702
rect 18604 29640 18656 29646
rect 18604 29582 18656 29588
rect 18696 29640 18748 29646
rect 19064 29640 19116 29646
rect 18748 29588 18828 29594
rect 18696 29582 18828 29588
rect 19064 29582 19116 29588
rect 18616 29306 18644 29582
rect 18708 29566 18828 29582
rect 19352 29578 19380 30144
rect 19536 29850 19564 30262
rect 19628 30190 19656 30330
rect 19892 30252 19944 30258
rect 19944 30212 20024 30240
rect 19892 30194 19944 30200
rect 19616 30184 19668 30190
rect 19616 30126 19668 30132
rect 19800 30116 19852 30122
rect 19800 30058 19852 30064
rect 19812 29850 19840 30058
rect 19524 29844 19576 29850
rect 19524 29786 19576 29792
rect 19800 29844 19852 29850
rect 19800 29786 19852 29792
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 18604 29300 18656 29306
rect 18604 29242 18656 29248
rect 18512 29232 18564 29238
rect 18512 29174 18564 29180
rect 18708 29170 18736 29446
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 18696 29164 18748 29170
rect 18696 29106 18748 29112
rect 17316 29028 17368 29034
rect 17316 28970 17368 28976
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 16580 27872 16632 27878
rect 16580 27814 16632 27820
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 16592 27538 16620 27814
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 17144 26994 17172 28018
rect 17328 27606 17356 28970
rect 17684 28076 17736 28082
rect 17684 28018 17736 28024
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17316 27600 17368 27606
rect 17316 27542 17368 27548
rect 17604 27402 17632 27814
rect 17696 27606 17724 28018
rect 18420 28008 18472 28014
rect 18420 27950 18472 27956
rect 18432 27674 18460 27950
rect 18420 27668 18472 27674
rect 18420 27610 18472 27616
rect 18800 27606 18828 29566
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 17684 27600 17736 27606
rect 17684 27542 17736 27548
rect 18788 27600 18840 27606
rect 18788 27542 18840 27548
rect 17960 27532 18012 27538
rect 17960 27474 18012 27480
rect 17684 27464 17736 27470
rect 17684 27406 17736 27412
rect 17776 27464 17828 27470
rect 17776 27406 17828 27412
rect 17592 27396 17644 27402
rect 17592 27338 17644 27344
rect 17132 26988 17184 26994
rect 17132 26930 17184 26936
rect 17500 26920 17552 26926
rect 17604 26908 17632 27338
rect 17552 26880 17632 26908
rect 17696 26908 17724 27406
rect 17788 27130 17816 27406
rect 17776 27124 17828 27130
rect 17776 27066 17828 27072
rect 17972 26994 18000 27474
rect 18328 27396 18380 27402
rect 18328 27338 18380 27344
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 17776 26920 17828 26926
rect 17696 26880 17776 26908
rect 17500 26862 17552 26868
rect 17776 26862 17828 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 16304 24812 16356 24818
rect 16304 24754 16356 24760
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 16316 24410 16344 24754
rect 16304 24404 16356 24410
rect 16304 24346 16356 24352
rect 16960 24206 16988 25842
rect 17236 25498 17264 26250
rect 17512 25838 17540 26862
rect 17788 26314 17816 26862
rect 17972 26382 18000 26930
rect 18340 26586 18368 27338
rect 18512 27328 18564 27334
rect 18512 27270 18564 27276
rect 18524 26994 18552 27270
rect 18512 26988 18564 26994
rect 18512 26930 18564 26936
rect 18512 26784 18564 26790
rect 18512 26726 18564 26732
rect 18328 26580 18380 26586
rect 18328 26522 18380 26528
rect 18236 26444 18288 26450
rect 18236 26386 18288 26392
rect 17960 26376 18012 26382
rect 17960 26318 18012 26324
rect 17776 26308 17828 26314
rect 17776 26250 17828 26256
rect 17500 25832 17552 25838
rect 17500 25774 17552 25780
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17316 25356 17368 25362
rect 17316 25298 17368 25304
rect 17040 24676 17092 24682
rect 17040 24618 17092 24624
rect 17052 24562 17080 24618
rect 17328 24614 17356 25298
rect 17408 25288 17460 25294
rect 17408 25230 17460 25236
rect 17420 24886 17448 25230
rect 17408 24880 17460 24886
rect 17408 24822 17460 24828
rect 17316 24608 17368 24614
rect 17052 24534 17264 24562
rect 17316 24550 17368 24556
rect 17236 24274 17264 24534
rect 17328 24342 17356 24550
rect 17316 24336 17368 24342
rect 17316 24278 17368 24284
rect 17512 24274 17540 25774
rect 17960 25764 18012 25770
rect 17960 25706 18012 25712
rect 17972 25362 18000 25706
rect 17960 25356 18012 25362
rect 17960 25298 18012 25304
rect 18248 25294 18276 26386
rect 18524 26382 18552 26726
rect 18800 26450 18828 27542
rect 19260 26994 19288 29174
rect 19352 29170 19380 29514
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19340 29164 19392 29170
rect 19340 29106 19392 29112
rect 19352 27878 19380 29106
rect 19996 29102 20024 30212
rect 20088 30054 20116 31282
rect 20260 31136 20312 31142
rect 20260 31078 20312 31084
rect 20272 30734 20300 31078
rect 20352 30932 20404 30938
rect 20352 30874 20404 30880
rect 20260 30728 20312 30734
rect 20260 30670 20312 30676
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20076 30048 20128 30054
rect 20076 29990 20128 29996
rect 20180 29782 20208 30602
rect 20272 30394 20300 30670
rect 20364 30598 20392 30874
rect 21376 30734 21404 31826
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22836 31272 22888 31278
rect 22836 31214 22888 31220
rect 21732 31136 21784 31142
rect 21732 31078 21784 31084
rect 22376 31136 22428 31142
rect 22376 31078 22428 31084
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21744 30666 21772 31078
rect 22008 30728 22060 30734
rect 22008 30670 22060 30676
rect 21732 30660 21784 30666
rect 21732 30602 21784 30608
rect 20352 30592 20404 30598
rect 20352 30534 20404 30540
rect 20260 30388 20312 30394
rect 20260 30330 20312 30336
rect 20364 29850 20392 30534
rect 22020 30326 22048 30670
rect 22008 30320 22060 30326
rect 22008 30262 22060 30268
rect 21916 30184 21968 30190
rect 21916 30126 21968 30132
rect 20812 30116 20864 30122
rect 20812 30058 20864 30064
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20168 29776 20220 29782
rect 20168 29718 20220 29724
rect 20824 29714 20852 30058
rect 21088 30048 21140 30054
rect 21088 29990 21140 29996
rect 20812 29708 20864 29714
rect 20812 29650 20864 29656
rect 21100 29646 21128 29990
rect 21928 29782 21956 30126
rect 21456 29776 21508 29782
rect 21456 29718 21508 29724
rect 21916 29776 21968 29782
rect 21916 29718 21968 29724
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20088 29238 20116 29582
rect 20168 29572 20220 29578
rect 20168 29514 20220 29520
rect 20180 29306 20208 29514
rect 20168 29300 20220 29306
rect 20168 29242 20220 29248
rect 20076 29232 20128 29238
rect 20076 29174 20128 29180
rect 19984 29096 20036 29102
rect 19984 29038 20036 29044
rect 19892 28552 19944 28558
rect 19996 28540 20024 29038
rect 19944 28512 20024 28540
rect 19892 28494 19944 28500
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19340 27872 19392 27878
rect 19340 27814 19392 27820
rect 19064 26988 19116 26994
rect 19064 26930 19116 26936
rect 19248 26988 19300 26994
rect 19248 26930 19300 26936
rect 19076 26586 19104 26930
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 18788 26444 18840 26450
rect 18788 26386 18840 26392
rect 18512 26376 18564 26382
rect 18512 26318 18564 26324
rect 19260 26314 19288 26930
rect 19352 26858 19380 27814
rect 19996 27470 20024 28512
rect 20168 28484 20220 28490
rect 20168 28426 20220 28432
rect 20180 28150 20208 28426
rect 21180 28416 21232 28422
rect 21180 28358 21232 28364
rect 20168 28144 20220 28150
rect 20168 28086 20220 28092
rect 21192 28082 21220 28358
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 21180 28076 21232 28082
rect 21180 28018 21232 28024
rect 20640 27606 20668 28018
rect 21468 28014 21496 29718
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21836 28994 21864 29650
rect 22020 29102 22048 30262
rect 22192 30184 22244 30190
rect 22192 30126 22244 30132
rect 22204 29850 22232 30126
rect 22192 29844 22244 29850
rect 22192 29786 22244 29792
rect 22100 29572 22152 29578
rect 22100 29514 22152 29520
rect 22008 29096 22060 29102
rect 22008 29038 22060 29044
rect 21836 28966 21956 28994
rect 21928 28626 21956 28966
rect 21916 28620 21968 28626
rect 21916 28562 21968 28568
rect 21824 28552 21876 28558
rect 22112 28540 22140 29514
rect 22388 29510 22416 31078
rect 22848 30938 22876 31214
rect 22468 30932 22520 30938
rect 22468 30874 22520 30880
rect 22836 30932 22888 30938
rect 22836 30874 22888 30880
rect 22480 30258 22508 30874
rect 22848 30258 22876 30874
rect 22468 30252 22520 30258
rect 22468 30194 22520 30200
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22480 29646 22508 30194
rect 22848 29646 22876 30194
rect 22940 29850 22968 31282
rect 23480 30184 23532 30190
rect 23480 30126 23532 30132
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 22468 29640 22520 29646
rect 22468 29582 22520 29588
rect 22836 29640 22888 29646
rect 22836 29582 22888 29588
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23216 29510 23244 29582
rect 23492 29578 23520 30126
rect 24228 29646 24256 32234
rect 24400 32224 24452 32230
rect 24400 32166 24452 32172
rect 24216 29640 24268 29646
rect 24216 29582 24268 29588
rect 23480 29572 23532 29578
rect 23480 29514 23532 29520
rect 22284 29504 22336 29510
rect 22284 29446 22336 29452
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 23204 29504 23256 29510
rect 23204 29446 23256 29452
rect 22296 28762 22324 29446
rect 22388 29170 22416 29446
rect 22376 29164 22428 29170
rect 22376 29106 22428 29112
rect 23216 28762 23244 29446
rect 22284 28756 22336 28762
rect 22284 28698 22336 28704
rect 22652 28756 22704 28762
rect 22652 28698 22704 28704
rect 23204 28756 23256 28762
rect 23204 28698 23256 28704
rect 22192 28552 22244 28558
rect 22112 28512 22192 28540
rect 21824 28494 21876 28500
rect 22192 28494 22244 28500
rect 21836 28422 21864 28494
rect 22664 28490 22692 28698
rect 22744 28688 22796 28694
rect 22744 28630 22796 28636
rect 22652 28484 22704 28490
rect 22652 28426 22704 28432
rect 21824 28416 21876 28422
rect 21824 28358 21876 28364
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 21456 28008 21508 28014
rect 21456 27950 21508 27956
rect 22112 27946 22140 28358
rect 22664 28014 22692 28426
rect 22652 28008 22704 28014
rect 22652 27950 22704 27956
rect 22100 27940 22152 27946
rect 22100 27882 22152 27888
rect 22560 27940 22612 27946
rect 22560 27882 22612 27888
rect 22284 27872 22336 27878
rect 22284 27814 22336 27820
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 22296 27470 22324 27814
rect 19984 27464 20036 27470
rect 19984 27406 20036 27412
rect 22284 27464 22336 27470
rect 22284 27406 22336 27412
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19340 26852 19392 26858
rect 19340 26794 19392 26800
rect 19248 26308 19300 26314
rect 19248 26250 19300 26256
rect 19352 25974 19380 26794
rect 19996 26790 20024 27406
rect 22572 26994 22600 27882
rect 22664 27674 22692 27950
rect 22652 27668 22704 27674
rect 22652 27610 22704 27616
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22100 26920 22152 26926
rect 22100 26862 22152 26868
rect 21364 26852 21416 26858
rect 21364 26794 21416 26800
rect 19984 26784 20036 26790
rect 19984 26726 20036 26732
rect 21088 26784 21140 26790
rect 21088 26726 21140 26732
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19340 25968 19392 25974
rect 19392 25928 19472 25956
rect 19340 25910 19392 25916
rect 19340 25832 19392 25838
rect 19340 25774 19392 25780
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 17684 25288 17736 25294
rect 17684 25230 17736 25236
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18788 25288 18840 25294
rect 18788 25230 18840 25236
rect 17696 24410 17724 25230
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 17868 24880 17920 24886
rect 17868 24822 17920 24828
rect 17776 24812 17828 24818
rect 17776 24754 17828 24760
rect 17684 24404 17736 24410
rect 17684 24346 17736 24352
rect 17224 24268 17276 24274
rect 17224 24210 17276 24216
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 16948 24200 17000 24206
rect 16948 24142 17000 24148
rect 17236 23866 17264 24210
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 17788 23798 17816 24754
rect 17880 24206 17908 24822
rect 18616 24818 18644 25094
rect 18800 24818 18828 25230
rect 19076 24818 19104 25298
rect 19248 25220 19300 25226
rect 19248 25162 19300 25168
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18788 24812 18840 24818
rect 18788 24754 18840 24760
rect 19064 24812 19116 24818
rect 19064 24754 19116 24760
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18708 24206 18736 24686
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 19260 24562 19288 25162
rect 19352 24682 19380 25774
rect 19340 24676 19392 24682
rect 19340 24618 19392 24624
rect 18800 24206 18828 24550
rect 19260 24534 19380 24562
rect 17868 24200 17920 24206
rect 17868 24142 17920 24148
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18788 24200 18840 24206
rect 18788 24142 18840 24148
rect 17776 23792 17828 23798
rect 17776 23734 17828 23740
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 17788 23118 17816 23734
rect 17776 23112 17828 23118
rect 17776 23054 17828 23060
rect 17880 22778 17908 24142
rect 18236 24064 18288 24070
rect 18236 24006 18288 24012
rect 18248 23730 18276 24006
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 19352 23118 19380 24534
rect 19444 24274 19472 25928
rect 19708 25900 19760 25906
rect 19708 25842 19760 25848
rect 19720 25498 19748 25842
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19892 25288 19944 25294
rect 19996 25242 20024 26726
rect 21100 26382 21128 26726
rect 21376 26586 21404 26794
rect 21364 26580 21416 26586
rect 21364 26522 21416 26528
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 20076 26308 20128 26314
rect 20076 26250 20128 26256
rect 20088 25906 20116 26250
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25786 20116 25842
rect 20088 25758 20300 25786
rect 20076 25696 20128 25702
rect 20076 25638 20128 25644
rect 20088 25294 20116 25638
rect 19944 25236 20024 25242
rect 19892 25230 20024 25236
rect 20076 25288 20128 25294
rect 20076 25230 20128 25236
rect 19904 25214 20024 25230
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19996 24818 20024 25214
rect 19984 24812 20036 24818
rect 19984 24754 20036 24760
rect 20168 24812 20220 24818
rect 20168 24754 20220 24760
rect 20180 24410 20208 24754
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 19432 24268 19484 24274
rect 19432 24210 19484 24216
rect 19444 23730 19472 24210
rect 20272 24206 20300 25758
rect 21376 25226 21404 26522
rect 22112 25498 22140 26862
rect 22204 25974 22232 26930
rect 22664 26926 22692 27610
rect 22756 27130 22784 28630
rect 23112 28552 23164 28558
rect 23112 28494 23164 28500
rect 23124 28150 23152 28494
rect 23112 28144 23164 28150
rect 23112 28086 23164 28092
rect 23124 27878 23152 28086
rect 23112 27872 23164 27878
rect 23112 27814 23164 27820
rect 22744 27124 22796 27130
rect 22744 27066 22796 27072
rect 22652 26920 22704 26926
rect 22652 26862 22704 26868
rect 23124 26382 23152 27814
rect 23492 27538 23520 29514
rect 23756 29300 23808 29306
rect 23756 29242 23808 29248
rect 23572 28960 23624 28966
rect 23572 28902 23624 28908
rect 23584 28558 23612 28902
rect 23768 28762 23796 29242
rect 24412 28762 24440 32166
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 24400 28756 24452 28762
rect 24400 28698 24452 28704
rect 23572 28552 23624 28558
rect 23572 28494 23624 28500
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23676 28218 23704 28494
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23584 27606 23612 27950
rect 23572 27600 23624 27606
rect 23572 27542 23624 27548
rect 23480 27532 23532 27538
rect 23480 27474 23532 27480
rect 23676 27470 23704 28154
rect 24412 28014 24440 28698
rect 24504 28082 24532 37062
rect 32324 36922 32352 37198
rect 32312 36916 32364 36922
rect 32312 36858 32364 36864
rect 32496 36780 32548 36786
rect 32496 36722 32548 36728
rect 32508 35894 32536 36722
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 32324 35866 32536 35894
rect 26976 34128 27028 34134
rect 26976 34070 27028 34076
rect 31208 34128 31260 34134
rect 31208 34070 31260 34076
rect 26792 34060 26844 34066
rect 26792 34002 26844 34008
rect 25136 33992 25188 33998
rect 25136 33934 25188 33940
rect 26516 33992 26568 33998
rect 26516 33934 26568 33940
rect 24860 33924 24912 33930
rect 24860 33866 24912 33872
rect 24872 33522 24900 33866
rect 24860 33516 24912 33522
rect 24860 33458 24912 33464
rect 24872 33046 24900 33458
rect 25148 33386 25176 33934
rect 26528 33658 26556 33934
rect 26516 33652 26568 33658
rect 26516 33594 26568 33600
rect 26056 33448 26108 33454
rect 26056 33390 26108 33396
rect 25136 33380 25188 33386
rect 25136 33322 25188 33328
rect 24860 33040 24912 33046
rect 24860 32982 24912 32988
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 24596 30734 24624 32914
rect 25148 32910 25176 33322
rect 24860 32904 24912 32910
rect 24860 32846 24912 32852
rect 25136 32904 25188 32910
rect 25136 32846 25188 32852
rect 25228 32904 25280 32910
rect 25228 32846 25280 32852
rect 25964 32904 26016 32910
rect 25964 32846 26016 32852
rect 24872 32298 24900 32846
rect 25044 32836 25096 32842
rect 25044 32778 25096 32784
rect 24952 32768 25004 32774
rect 24952 32710 25004 32716
rect 24860 32292 24912 32298
rect 24860 32234 24912 32240
rect 24768 32224 24820 32230
rect 24768 32166 24820 32172
rect 24780 31958 24808 32166
rect 24768 31952 24820 31958
rect 24768 31894 24820 31900
rect 24964 30938 24992 32710
rect 25056 31822 25084 32778
rect 25240 32570 25268 32846
rect 25976 32570 26004 32846
rect 26068 32722 26096 33390
rect 26528 33318 26556 33594
rect 26516 33312 26568 33318
rect 26516 33254 26568 33260
rect 26528 32774 26556 33254
rect 26804 33114 26832 34002
rect 26792 33108 26844 33114
rect 26792 33050 26844 33056
rect 26988 32910 27016 34070
rect 27620 33992 27672 33998
rect 27620 33934 27672 33940
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28540 33992 28592 33998
rect 28540 33934 28592 33940
rect 29184 33992 29236 33998
rect 29184 33934 29236 33940
rect 30104 33992 30156 33998
rect 30104 33934 30156 33940
rect 31024 33992 31076 33998
rect 31024 33934 31076 33940
rect 27632 33658 27660 33934
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27252 33516 27304 33522
rect 27252 33458 27304 33464
rect 27620 33516 27672 33522
rect 27620 33458 27672 33464
rect 27264 32910 27292 33458
rect 27632 33114 27660 33458
rect 27620 33108 27672 33114
rect 27620 33050 27672 33056
rect 28276 32978 28304 33934
rect 28356 33856 28408 33862
rect 28356 33798 28408 33804
rect 28448 33856 28500 33862
rect 28448 33798 28500 33804
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 27252 32904 27304 32910
rect 27252 32846 27304 32852
rect 26516 32768 26568 32774
rect 26068 32694 26188 32722
rect 26516 32710 26568 32716
rect 25228 32564 25280 32570
rect 25228 32506 25280 32512
rect 25964 32564 26016 32570
rect 25964 32506 26016 32512
rect 25136 32428 25188 32434
rect 25136 32370 25188 32376
rect 25780 32428 25832 32434
rect 25780 32370 25832 32376
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 24952 30932 25004 30938
rect 24952 30874 25004 30880
rect 24584 30728 24636 30734
rect 24584 30670 24636 30676
rect 25044 30728 25096 30734
rect 25148 30716 25176 32370
rect 25228 32292 25280 32298
rect 25228 32234 25280 32240
rect 25240 31822 25268 32234
rect 25792 32230 25820 32370
rect 26160 32366 26188 32694
rect 26148 32360 26200 32366
rect 26148 32302 26200 32308
rect 25780 32224 25832 32230
rect 25780 32166 25832 32172
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 26056 31816 26108 31822
rect 26056 31758 26108 31764
rect 26160 31770 26188 32302
rect 27264 31958 27292 32846
rect 28172 32428 28224 32434
rect 28172 32370 28224 32376
rect 27620 32360 27672 32366
rect 27620 32302 27672 32308
rect 27252 31952 27304 31958
rect 26344 31878 26556 31906
rect 27252 31894 27304 31900
rect 27436 31952 27488 31958
rect 27436 31894 27488 31900
rect 26344 31770 26372 31878
rect 26068 31346 26096 31758
rect 26160 31742 26372 31770
rect 26528 31754 26556 31878
rect 27448 31754 27476 31894
rect 27632 31754 27660 32302
rect 28080 32224 28132 32230
rect 28080 32166 28132 32172
rect 26528 31748 26660 31754
rect 26528 31726 26608 31748
rect 26608 31690 26660 31696
rect 27356 31726 27476 31754
rect 27620 31748 27672 31754
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26252 31482 26280 31622
rect 26240 31476 26292 31482
rect 26240 31418 26292 31424
rect 26056 31340 26108 31346
rect 26056 31282 26108 31288
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 25504 30932 25556 30938
rect 25504 30874 25556 30880
rect 25096 30688 25176 30716
rect 25044 30670 25096 30676
rect 24860 30592 24912 30598
rect 24860 30534 24912 30540
rect 24872 29850 24900 30534
rect 24952 30252 25004 30258
rect 24952 30194 25004 30200
rect 24964 29850 24992 30194
rect 25056 30054 25084 30670
rect 25516 30190 25544 30874
rect 25780 30796 25832 30802
rect 25780 30738 25832 30744
rect 25792 30190 25820 30738
rect 26240 30728 26292 30734
rect 26240 30670 26292 30676
rect 26608 30728 26660 30734
rect 26608 30670 26660 30676
rect 26884 30728 26936 30734
rect 26884 30670 26936 30676
rect 25872 30660 25924 30666
rect 25872 30602 25924 30608
rect 25504 30184 25556 30190
rect 25504 30126 25556 30132
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 24860 29844 24912 29850
rect 24860 29786 24912 29792
rect 24952 29844 25004 29850
rect 24952 29786 25004 29792
rect 24952 29708 25004 29714
rect 24952 29650 25004 29656
rect 24860 28620 24912 28626
rect 24860 28562 24912 28568
rect 24492 28076 24544 28082
rect 24492 28018 24544 28024
rect 24124 28008 24176 28014
rect 24124 27950 24176 27956
rect 24400 28008 24452 28014
rect 24400 27950 24452 27956
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23112 26376 23164 26382
rect 23112 26318 23164 26324
rect 22928 26240 22980 26246
rect 22928 26182 22980 26188
rect 22192 25968 22244 25974
rect 22192 25910 22244 25916
rect 22560 25968 22612 25974
rect 22560 25910 22612 25916
rect 22572 25498 22600 25910
rect 22100 25492 22152 25498
rect 22100 25434 22152 25440
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22468 25424 22520 25430
rect 22468 25366 22520 25372
rect 21916 25356 21968 25362
rect 21916 25298 21968 25304
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21928 25242 21956 25298
rect 21364 25220 21416 25226
rect 21364 25162 21416 25168
rect 21836 24750 21864 25230
rect 21928 25214 22048 25242
rect 22020 25158 22048 25214
rect 22008 25152 22060 25158
rect 22008 25094 22060 25100
rect 22284 25152 22336 25158
rect 22284 25094 22336 25100
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 21824 24744 21876 24750
rect 21824 24686 21876 24692
rect 21272 24608 21324 24614
rect 21272 24550 21324 24556
rect 21284 24206 21312 24550
rect 22020 24206 22048 24890
rect 22100 24812 22152 24818
rect 22100 24754 22152 24760
rect 22112 24206 22140 24754
rect 22296 24410 22324 25094
rect 22480 24818 22508 25366
rect 22940 25294 22968 26182
rect 23124 26042 23152 26318
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 23112 25900 23164 25906
rect 23112 25842 23164 25848
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22928 25288 22980 25294
rect 22928 25230 22980 25236
rect 22468 24812 22520 24818
rect 22468 24754 22520 24760
rect 22664 24682 22692 25230
rect 23124 25226 23152 25842
rect 23204 25696 23256 25702
rect 23204 25638 23256 25644
rect 23216 25294 23244 25638
rect 23204 25288 23256 25294
rect 23204 25230 23256 25236
rect 23112 25220 23164 25226
rect 23112 25162 23164 25168
rect 22652 24676 22704 24682
rect 22652 24618 22704 24624
rect 22284 24404 22336 24410
rect 22284 24346 22336 24352
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 19984 24200 20036 24206
rect 20260 24200 20312 24206
rect 19984 24142 20036 24148
rect 20258 24168 20260 24177
rect 21272 24200 21324 24206
rect 20312 24168 20314 24177
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19996 23866 20024 24142
rect 21272 24142 21324 24148
rect 21640 24200 21692 24206
rect 21640 24142 21692 24148
rect 22008 24200 22060 24206
rect 22008 24142 22060 24148
rect 22100 24200 22152 24206
rect 22100 24142 22152 24148
rect 20258 24103 20314 24112
rect 19984 23860 20036 23866
rect 19984 23802 20036 23808
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19444 23322 19472 23666
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 18604 23044 18656 23050
rect 18604 22986 18656 22992
rect 17960 22976 18012 22982
rect 17960 22918 18012 22924
rect 17868 22772 17920 22778
rect 17868 22714 17920 22720
rect 17972 22642 18000 22918
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17880 21554 17908 22034
rect 17972 22030 18000 22578
rect 17960 22024 18012 22030
rect 17960 21966 18012 21972
rect 18064 21894 18092 22714
rect 18616 22642 18644 22986
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 19340 22976 19392 22982
rect 19340 22918 19392 22924
rect 18800 22778 18828 22918
rect 18788 22772 18840 22778
rect 18788 22714 18840 22720
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18604 22636 18656 22642
rect 18604 22578 18656 22584
rect 18156 21962 18184 22578
rect 18800 22234 18828 22714
rect 19352 22658 19380 22918
rect 19444 22778 19472 23258
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19432 22772 19484 22778
rect 19432 22714 19484 22720
rect 19168 22642 19380 22658
rect 19156 22636 19380 22642
rect 19208 22630 19380 22636
rect 19156 22578 19208 22584
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 19432 22568 19484 22574
rect 19432 22510 19484 22516
rect 18788 22228 18840 22234
rect 18788 22170 18840 22176
rect 18144 21956 18196 21962
rect 18144 21898 18196 21904
rect 18052 21888 18104 21894
rect 18880 21888 18932 21894
rect 18052 21830 18104 21836
rect 18800 21848 18880 21876
rect 18800 21554 18828 21848
rect 18880 21830 18932 21836
rect 19076 21690 19104 22510
rect 19064 21684 19116 21690
rect 19064 21626 19116 21632
rect 19444 21554 19472 22510
rect 19996 22438 20024 23054
rect 20272 22982 20300 24103
rect 21652 23866 21680 24142
rect 22204 24126 22508 24154
rect 21640 23860 21692 23866
rect 21640 23802 21692 23808
rect 22204 23730 22232 24126
rect 22480 24070 22508 24126
rect 22376 24064 22428 24070
rect 22376 24006 22428 24012
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22388 23730 22416 24006
rect 22572 23730 22600 24210
rect 21272 23724 21324 23730
rect 21272 23666 21324 23672
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 22192 23724 22244 23730
rect 22192 23666 22244 23672
rect 22376 23724 22428 23730
rect 22376 23666 22428 23672
rect 22560 23724 22612 23730
rect 22560 23666 22612 23672
rect 20444 23316 20496 23322
rect 20444 23258 20496 23264
rect 20260 22976 20312 22982
rect 20260 22918 20312 22924
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21570 20024 22374
rect 20456 22234 20484 23258
rect 20812 23180 20864 23186
rect 20812 23122 20864 23128
rect 20720 23112 20772 23118
rect 20824 23089 20852 23122
rect 20720 23054 20772 23060
rect 20810 23080 20866 23089
rect 20444 22228 20496 22234
rect 20444 22170 20496 22176
rect 20732 22030 20760 23054
rect 21284 23050 21312 23666
rect 21824 23656 21876 23662
rect 21652 23604 21824 23610
rect 21652 23598 21876 23604
rect 21652 23582 21864 23598
rect 21652 23526 21680 23582
rect 21640 23520 21692 23526
rect 21640 23462 21692 23468
rect 21652 23118 21680 23462
rect 22020 23322 22048 23666
rect 22008 23316 22060 23322
rect 22008 23258 22060 23264
rect 21640 23112 21692 23118
rect 21640 23054 21692 23060
rect 21824 23112 21876 23118
rect 21916 23112 21968 23118
rect 21824 23054 21876 23060
rect 21914 23080 21916 23089
rect 21968 23080 21970 23089
rect 20810 23015 20866 23024
rect 21272 23044 21324 23050
rect 21272 22986 21324 22992
rect 21284 22778 21312 22986
rect 21364 22976 21416 22982
rect 21364 22918 21416 22924
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21376 22438 21404 22918
rect 21836 22778 21864 23054
rect 22204 23050 22232 23666
rect 21914 23015 21970 23024
rect 22192 23044 22244 23050
rect 22192 22986 22244 22992
rect 21824 22772 21876 22778
rect 21824 22714 21876 22720
rect 22204 22438 22232 22986
rect 22388 22710 22416 23666
rect 22664 23594 22692 24618
rect 23124 24206 23152 25162
rect 23216 24274 23244 25230
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23112 24200 23164 24206
rect 23112 24142 23164 24148
rect 22652 23588 22704 23594
rect 22652 23530 22704 23536
rect 22664 23186 22692 23530
rect 22652 23180 22704 23186
rect 22652 23122 22704 23128
rect 22928 23044 22980 23050
rect 22928 22986 22980 22992
rect 22940 22778 22968 22986
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22376 22704 22428 22710
rect 22376 22646 22428 22652
rect 23124 22642 23152 24142
rect 23400 23798 23428 25842
rect 23756 24336 23808 24342
rect 23756 24278 23808 24284
rect 23572 24268 23624 24274
rect 23572 24210 23624 24216
rect 23388 23792 23440 23798
rect 23388 23734 23440 23740
rect 23112 22636 23164 22642
rect 23112 22578 23164 22584
rect 23124 22506 23152 22578
rect 23112 22500 23164 22506
rect 23112 22442 23164 22448
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 22192 22432 22244 22438
rect 22192 22374 22244 22380
rect 22560 22432 22612 22438
rect 22560 22374 22612 22380
rect 21376 22030 21404 22374
rect 22572 22030 22600 22374
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 21364 22024 21416 22030
rect 21364 21966 21416 21972
rect 22560 22024 22612 22030
rect 22560 21966 22612 21972
rect 23112 22024 23164 22030
rect 23164 21972 23244 21978
rect 23112 21966 23244 21972
rect 20904 21956 20956 21962
rect 20904 21898 20956 21904
rect 20076 21888 20128 21894
rect 20076 21830 20128 21836
rect 19904 21554 20024 21570
rect 20088 21554 20116 21830
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 18788 21548 18840 21554
rect 18788 21490 18840 21496
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19892 21548 20024 21554
rect 19944 21542 20024 21548
rect 20076 21548 20128 21554
rect 19892 21490 19944 21496
rect 20076 21490 20128 21496
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 1768 20936 1820 20942
rect 1768 20878 1820 20884
rect 1780 20505 1808 20878
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 1766 20496 1822 20505
rect 1766 20431 1822 20440
rect 20628 20460 20680 20466
rect 20628 20402 20680 20408
rect 20076 20256 20128 20262
rect 20076 20198 20128 20204
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 19432 19848 19484 19854
rect 19432 19790 19484 19796
rect 19444 19446 19472 19790
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19432 19440 19484 19446
rect 19432 19382 19484 19388
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 19444 18766 19472 19382
rect 19708 19168 19760 19174
rect 19708 19110 19760 19116
rect 19720 18766 19748 19110
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19708 18760 19760 18766
rect 19708 18702 19760 18708
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 19444 17202 19472 18702
rect 19984 18692 20036 18698
rect 19984 18634 20036 18640
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19996 18290 20024 18634
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19984 17536 20036 17542
rect 19984 17478 20036 17484
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19996 17270 20024 17478
rect 19984 17264 20036 17270
rect 19984 17206 20036 17212
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 20088 16114 20116 20198
rect 20352 19780 20404 19786
rect 20352 19722 20404 19728
rect 20364 19514 20392 19722
rect 20352 19508 20404 19514
rect 20352 19450 20404 19456
rect 20548 19378 20576 20198
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20180 18426 20208 19246
rect 20640 18698 20668 20402
rect 20720 19304 20772 19310
rect 20720 19246 20772 19252
rect 20628 18692 20680 18698
rect 20628 18634 20680 18640
rect 20168 18420 20220 18426
rect 20168 18362 20220 18368
rect 20732 18154 20760 19246
rect 20812 19168 20864 19174
rect 20812 19110 20864 19116
rect 20824 18426 20852 19110
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20720 18148 20772 18154
rect 20720 18090 20772 18096
rect 20732 17882 20760 18090
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20732 17678 20760 17818
rect 20444 17672 20496 17678
rect 20444 17614 20496 17620
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 20456 17542 20484 17614
rect 20916 17610 20944 21898
rect 21192 21690 21220 21966
rect 23124 21950 23244 21966
rect 23216 21894 23244 21950
rect 22100 21888 22152 21894
rect 22100 21830 22152 21836
rect 23204 21888 23256 21894
rect 23204 21830 23256 21836
rect 21180 21684 21232 21690
rect 21180 21626 21232 21632
rect 22112 21622 22140 21830
rect 23216 21690 23244 21830
rect 23204 21684 23256 21690
rect 23204 21626 23256 21632
rect 22100 21616 22152 21622
rect 22100 21558 22152 21564
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 22020 20942 22048 21490
rect 22008 20936 22060 20942
rect 22008 20878 22060 20884
rect 22192 19848 22244 19854
rect 22192 19790 22244 19796
rect 21640 19780 21692 19786
rect 21640 19722 21692 19728
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19310 21312 19654
rect 21272 19304 21324 19310
rect 21272 19246 21324 19252
rect 21284 18766 21312 19246
rect 21652 19174 21680 19722
rect 22008 19372 22060 19378
rect 22008 19314 22060 19320
rect 21640 19168 21692 19174
rect 21640 19110 21692 19116
rect 21652 18766 21680 19110
rect 22020 18766 22048 19314
rect 21272 18760 21324 18766
rect 21272 18702 21324 18708
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 22008 18760 22060 18766
rect 22008 18702 22060 18708
rect 21180 18624 21232 18630
rect 21180 18566 21232 18572
rect 21192 18358 21220 18566
rect 21180 18352 21232 18358
rect 21180 18294 21232 18300
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20444 17536 20496 17542
rect 20444 17478 20496 17484
rect 20456 16998 20484 17478
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20444 16992 20496 16998
rect 20444 16934 20496 16940
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20180 16182 20208 16934
rect 20640 16726 20668 16934
rect 20444 16720 20496 16726
rect 20444 16662 20496 16668
rect 20628 16720 20680 16726
rect 20628 16662 20680 16668
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20168 16176 20220 16182
rect 20168 16118 20220 16124
rect 20076 16108 20128 16114
rect 20076 16050 20128 16056
rect 20272 15910 20300 16526
rect 20456 16046 20484 16662
rect 20720 16584 20772 16590
rect 20640 16544 20720 16572
rect 20640 16250 20668 16544
rect 20720 16526 20772 16532
rect 21192 16522 21220 18294
rect 21284 18086 21312 18702
rect 21272 18080 21324 18086
rect 21272 18022 21324 18028
rect 21284 16726 21312 18022
rect 21652 17814 21680 18702
rect 22204 18426 22232 19790
rect 22284 19712 22336 19718
rect 22284 19654 22336 19660
rect 22296 19446 22324 19654
rect 22284 19440 22336 19446
rect 22284 19382 22336 19388
rect 22376 19168 22428 19174
rect 22376 19110 22428 19116
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22388 18290 22416 19110
rect 23112 18624 23164 18630
rect 23112 18566 23164 18572
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22100 18216 22152 18222
rect 22100 18158 22152 18164
rect 21640 17808 21692 17814
rect 21640 17750 21692 17756
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21180 16516 21232 16522
rect 21180 16458 21232 16464
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 20628 16244 20680 16250
rect 20628 16186 20680 16192
rect 20444 16040 20496 16046
rect 20444 15982 20496 15988
rect 19340 15904 19392 15910
rect 19340 15846 19392 15852
rect 20260 15904 20312 15910
rect 20260 15846 20312 15852
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 1860 15700 1912 15706
rect 1860 15642 1912 15648
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1780 10305 1808 10406
rect 1766 10296 1822 10305
rect 1766 10231 1822 10240
rect 1872 2514 1900 15642
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 19352 6914 19380 15846
rect 20456 15706 20484 15982
rect 20444 15700 20496 15706
rect 20444 15642 20496 15648
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19444 14482 19472 14962
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 20088 13938 20116 14214
rect 20456 14074 20484 14282
rect 20444 14068 20496 14074
rect 20444 14010 20496 14016
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19892 13932 19944 13938
rect 19892 13874 19944 13880
rect 20076 13932 20128 13938
rect 20076 13874 20128 13880
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19444 12238 19472 13806
rect 19536 13462 19564 13874
rect 19800 13728 19852 13734
rect 19800 13670 19852 13676
rect 19524 13456 19576 13462
rect 19524 13398 19576 13404
rect 19812 13326 19840 13670
rect 19904 13530 19932 13874
rect 19892 13524 19944 13530
rect 19892 13466 19944 13472
rect 20456 13326 20484 13874
rect 20640 13530 20668 16186
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 20916 15706 20944 16050
rect 21008 15978 21036 16390
rect 21192 16114 21220 16458
rect 21284 16182 21312 16662
rect 21272 16176 21324 16182
rect 21272 16118 21324 16124
rect 22112 16114 22140 18158
rect 22388 17610 22416 18226
rect 23124 17678 23152 18566
rect 23400 18290 23428 23734
rect 23584 22710 23612 24210
rect 23572 22704 23624 22710
rect 23572 22646 23624 22652
rect 23584 22030 23612 22646
rect 23768 22642 23796 24278
rect 23848 24132 23900 24138
rect 23848 24074 23900 24080
rect 23860 23322 23888 24074
rect 23848 23316 23900 23322
rect 23848 23258 23900 23264
rect 24032 22704 24084 22710
rect 24032 22646 24084 22652
rect 23756 22636 23808 22642
rect 23756 22578 23808 22584
rect 23572 22024 23624 22030
rect 23572 21966 23624 21972
rect 23584 21554 23612 21966
rect 24044 21554 24072 22646
rect 23572 21548 23624 21554
rect 23572 21490 23624 21496
rect 24032 21548 24084 21554
rect 24032 21490 24084 21496
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 20874 23520 21286
rect 23584 21146 23612 21490
rect 23572 21140 23624 21146
rect 23572 21082 23624 21088
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23480 20868 23532 20874
rect 23480 20810 23532 20816
rect 23480 19712 23532 19718
rect 23480 19654 23532 19660
rect 23492 18698 23520 19654
rect 23584 18766 23612 20878
rect 24044 20534 24072 21490
rect 24032 20528 24084 20534
rect 24032 20470 24084 20476
rect 24044 20330 24072 20470
rect 24032 20324 24084 20330
rect 24032 20266 24084 20272
rect 23848 19848 23900 19854
rect 23848 19790 23900 19796
rect 24032 19848 24084 19854
rect 24032 19790 24084 19796
rect 23572 18760 23624 18766
rect 23572 18702 23624 18708
rect 23480 18692 23532 18698
rect 23480 18634 23532 18640
rect 23584 18426 23612 18702
rect 23572 18420 23624 18426
rect 23572 18362 23624 18368
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 22652 17672 22704 17678
rect 22652 17614 22704 17620
rect 23112 17672 23164 17678
rect 23112 17614 23164 17620
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 22192 17604 22244 17610
rect 22192 17546 22244 17552
rect 22376 17604 22428 17610
rect 22376 17546 22428 17552
rect 22204 16794 22232 17546
rect 22664 17202 22692 17614
rect 23308 17202 23336 17614
rect 23400 17270 23428 18226
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 22652 17196 22704 17202
rect 22652 17138 22704 17144
rect 23296 17196 23348 17202
rect 23296 17138 23348 17144
rect 22192 16788 22244 16794
rect 22192 16730 22244 16736
rect 22204 16590 22232 16730
rect 22192 16584 22244 16590
rect 22192 16526 22244 16532
rect 21180 16108 21232 16114
rect 21180 16050 21232 16056
rect 22100 16108 22152 16114
rect 22100 16050 22152 16056
rect 22376 16108 22428 16114
rect 22376 16050 22428 16056
rect 20996 15972 21048 15978
rect 20996 15914 21048 15920
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 22388 15638 22416 16050
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22664 15502 22692 17138
rect 23480 16720 23532 16726
rect 23480 16662 23532 16668
rect 22836 16584 22888 16590
rect 22836 16526 22888 16532
rect 22744 16448 22796 16454
rect 22744 16390 22796 16396
rect 22756 16250 22784 16390
rect 22744 16244 22796 16250
rect 22744 16186 22796 16192
rect 22848 15706 22876 16526
rect 23492 16522 23520 16662
rect 23112 16516 23164 16522
rect 23112 16458 23164 16464
rect 23480 16516 23532 16522
rect 23480 16458 23532 16464
rect 23124 15706 23152 16458
rect 23492 15706 23520 16458
rect 23584 16114 23612 18362
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23676 16658 23704 17478
rect 23860 17338 23888 19790
rect 24044 18086 24072 19790
rect 24136 18358 24164 27950
rect 24676 27328 24728 27334
rect 24676 27270 24728 27276
rect 24688 27062 24716 27270
rect 24676 27056 24728 27062
rect 24676 26998 24728 27004
rect 24676 26784 24728 26790
rect 24676 26726 24728 26732
rect 24688 26382 24716 26726
rect 24676 26376 24728 26382
rect 24676 26318 24728 26324
rect 24492 26308 24544 26314
rect 24492 26250 24544 26256
rect 24400 25832 24452 25838
rect 24400 25774 24452 25780
rect 24412 22710 24440 25774
rect 24504 25498 24532 26250
rect 24688 26042 24716 26318
rect 24676 26036 24728 26042
rect 24676 25978 24728 25984
rect 24492 25492 24544 25498
rect 24492 25434 24544 25440
rect 24584 25424 24636 25430
rect 24584 25366 24636 25372
rect 24492 25288 24544 25294
rect 24492 25230 24544 25236
rect 24504 24954 24532 25230
rect 24492 24948 24544 24954
rect 24492 24890 24544 24896
rect 24492 24812 24544 24818
rect 24492 24754 24544 24760
rect 24504 24410 24532 24754
rect 24492 24404 24544 24410
rect 24492 24346 24544 24352
rect 24596 24206 24624 25366
rect 24688 24886 24716 25978
rect 24872 25362 24900 28562
rect 24964 27470 24992 29650
rect 25056 29306 25084 29990
rect 25792 29646 25820 30126
rect 25884 29850 25912 30602
rect 26252 30326 26280 30670
rect 26240 30320 26292 30326
rect 26240 30262 26292 30268
rect 26620 30258 26648 30670
rect 26056 30252 26108 30258
rect 26056 30194 26108 30200
rect 26608 30252 26660 30258
rect 26608 30194 26660 30200
rect 26068 29850 26096 30194
rect 26896 30122 26924 30670
rect 27172 30258 27200 31282
rect 27252 30592 27304 30598
rect 27252 30534 27304 30540
rect 26976 30252 27028 30258
rect 26976 30194 27028 30200
rect 27160 30252 27212 30258
rect 27160 30194 27212 30200
rect 26884 30116 26936 30122
rect 26884 30058 26936 30064
rect 26988 30054 27016 30194
rect 26976 30048 27028 30054
rect 26976 29990 27028 29996
rect 25872 29844 25924 29850
rect 25872 29786 25924 29792
rect 26056 29844 26108 29850
rect 26056 29786 26108 29792
rect 26988 29646 27016 29990
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 26976 29640 27028 29646
rect 26976 29582 27028 29588
rect 25044 29300 25096 29306
rect 25044 29242 25096 29248
rect 25780 29164 25832 29170
rect 25780 29106 25832 29112
rect 26424 29164 26476 29170
rect 26424 29106 26476 29112
rect 25688 28960 25740 28966
rect 25688 28902 25740 28908
rect 25700 28490 25728 28902
rect 25688 28484 25740 28490
rect 25688 28426 25740 28432
rect 25792 28218 25820 29106
rect 26436 28762 26464 29106
rect 27068 29096 27120 29102
rect 27068 29038 27120 29044
rect 26424 28756 26476 28762
rect 26424 28698 26476 28704
rect 26240 28552 26292 28558
rect 26240 28494 26292 28500
rect 25780 28212 25832 28218
rect 25780 28154 25832 28160
rect 25044 28144 25096 28150
rect 25044 28086 25096 28092
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24964 25838 24992 27406
rect 24952 25832 25004 25838
rect 24952 25774 25004 25780
rect 24860 25356 24912 25362
rect 24860 25298 24912 25304
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24676 24880 24728 24886
rect 24676 24822 24728 24828
rect 24688 24274 24716 24822
rect 24676 24268 24728 24274
rect 24676 24210 24728 24216
rect 24780 24206 24808 25162
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24768 24200 24820 24206
rect 24768 24142 24820 24148
rect 24400 22704 24452 22710
rect 24400 22646 24452 22652
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24308 22568 24360 22574
rect 24308 22510 24360 22516
rect 24216 21548 24268 21554
rect 24216 21490 24268 21496
rect 24228 20466 24256 21490
rect 24320 21010 24348 22510
rect 24596 22234 24624 22578
rect 24584 22228 24636 22234
rect 24584 22170 24636 22176
rect 24872 22094 24900 25298
rect 24872 22066 24992 22094
rect 24308 21004 24360 21010
rect 24308 20946 24360 20952
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20602 24900 20810
rect 24860 20596 24912 20602
rect 24860 20538 24912 20544
rect 24216 20460 24268 20466
rect 24216 20402 24268 20408
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24216 19304 24268 19310
rect 24216 19246 24268 19252
rect 24228 18766 24256 19246
rect 24216 18760 24268 18766
rect 24216 18702 24268 18708
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24124 18352 24176 18358
rect 24124 18294 24176 18300
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17882 24072 18022
rect 24032 17876 24084 17882
rect 24032 17818 24084 17824
rect 24584 17672 24636 17678
rect 24584 17614 24636 17620
rect 23848 17332 23900 17338
rect 23848 17274 23900 17280
rect 24596 16794 24624 17614
rect 24688 17338 24716 18702
rect 24676 17332 24728 17338
rect 24676 17274 24728 17280
rect 24584 16788 24636 16794
rect 24584 16730 24636 16736
rect 24688 16658 24716 17274
rect 24872 17066 24900 20402
rect 24964 17134 24992 22066
rect 25056 21554 25084 28086
rect 25964 28076 26016 28082
rect 25964 28018 26016 28024
rect 25976 27878 26004 28018
rect 25964 27872 26016 27878
rect 25964 27814 26016 27820
rect 25688 27600 25740 27606
rect 25688 27542 25740 27548
rect 25228 27396 25280 27402
rect 25228 27338 25280 27344
rect 25240 21962 25268 27338
rect 25596 26308 25648 26314
rect 25596 26250 25648 26256
rect 25608 26042 25636 26250
rect 25596 26036 25648 26042
rect 25596 25978 25648 25984
rect 25700 25906 25728 27542
rect 26148 27396 26200 27402
rect 26148 27338 26200 27344
rect 26160 27062 26188 27338
rect 26148 27056 26200 27062
rect 26148 26998 26200 27004
rect 26160 26586 26188 26998
rect 26148 26580 26200 26586
rect 26148 26522 26200 26528
rect 26252 26382 26280 28494
rect 26436 28218 26464 28698
rect 27080 28218 27108 29038
rect 27172 28558 27200 30194
rect 27264 29646 27292 30534
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 27160 28552 27212 28558
rect 27160 28494 27212 28500
rect 27252 28552 27304 28558
rect 27252 28494 27304 28500
rect 26424 28212 26476 28218
rect 26424 28154 26476 28160
rect 27068 28212 27120 28218
rect 27068 28154 27120 28160
rect 26332 28076 26384 28082
rect 26332 28018 26384 28024
rect 26344 27470 26372 28018
rect 26332 27464 26384 27470
rect 26332 27406 26384 27412
rect 26344 27130 26372 27406
rect 26436 27334 26464 28154
rect 27264 27674 27292 28494
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27356 27538 27384 31726
rect 27620 31690 27672 31696
rect 27632 31482 27660 31690
rect 27620 31476 27672 31482
rect 27620 31418 27672 31424
rect 27632 30734 27660 31418
rect 28092 31414 28120 32166
rect 28080 31408 28132 31414
rect 28080 31350 28132 31356
rect 27620 30728 27672 30734
rect 27620 30670 27672 30676
rect 27436 30252 27488 30258
rect 27436 30194 27488 30200
rect 27448 29850 27476 30194
rect 27436 29844 27488 29850
rect 27436 29786 27488 29792
rect 27632 29578 27660 30670
rect 27620 29572 27672 29578
rect 27620 29514 27672 29520
rect 27620 29300 27672 29306
rect 27620 29242 27672 29248
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27344 27532 27396 27538
rect 27344 27474 27396 27480
rect 27448 27334 27476 28970
rect 27528 28416 27580 28422
rect 27528 28358 27580 28364
rect 27540 27470 27568 28358
rect 27528 27464 27580 27470
rect 27528 27406 27580 27412
rect 26424 27328 26476 27334
rect 26424 27270 26476 27276
rect 27436 27328 27488 27334
rect 27436 27270 27488 27276
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26436 26790 26464 27270
rect 27448 27130 27476 27270
rect 27436 27124 27488 27130
rect 27436 27066 27488 27072
rect 27632 26926 27660 29242
rect 27804 28960 27856 28966
rect 27804 28902 27856 28908
rect 27816 28490 27844 28902
rect 28080 28552 28132 28558
rect 28080 28494 28132 28500
rect 27804 28484 27856 28490
rect 27804 28426 27856 28432
rect 27896 28484 27948 28490
rect 27896 28426 27948 28432
rect 27908 28150 27936 28426
rect 27988 28416 28040 28422
rect 27988 28358 28040 28364
rect 27896 28144 27948 28150
rect 27896 28086 27948 28092
rect 28000 28082 28028 28358
rect 28092 28218 28120 28494
rect 28080 28212 28132 28218
rect 28080 28154 28132 28160
rect 27988 28076 28040 28082
rect 27988 28018 28040 28024
rect 28184 27470 28212 32370
rect 28368 31822 28396 33798
rect 28460 33454 28488 33798
rect 28448 33448 28500 33454
rect 28448 33390 28500 33396
rect 28552 32858 28580 33934
rect 29092 33380 29144 33386
rect 29092 33322 29144 33328
rect 28908 33312 28960 33318
rect 28908 33254 28960 33260
rect 28920 32978 28948 33254
rect 28908 32972 28960 32978
rect 28908 32914 28960 32920
rect 28460 32842 28580 32858
rect 28448 32836 28580 32842
rect 28500 32830 28580 32836
rect 28448 32778 28500 32784
rect 28460 32570 28488 32778
rect 28448 32564 28500 32570
rect 28448 32506 28500 32512
rect 28356 31816 28408 31822
rect 28356 31758 28408 31764
rect 28460 31142 28488 32506
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28540 32292 28592 32298
rect 28540 32234 28592 32240
rect 28448 31136 28500 31142
rect 28448 31078 28500 31084
rect 28460 29866 28488 31078
rect 28276 29838 28488 29866
rect 28276 29170 28304 29838
rect 28448 29640 28500 29646
rect 28448 29582 28500 29588
rect 28460 29510 28488 29582
rect 28448 29504 28500 29510
rect 28448 29446 28500 29452
rect 28552 29238 28580 32234
rect 28644 32230 28672 32370
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28644 31822 28672 32166
rect 28632 31816 28684 31822
rect 28632 31758 28684 31764
rect 28644 29782 28672 31758
rect 28920 31686 28948 32914
rect 29104 32434 29132 33322
rect 29196 33114 29224 33934
rect 30116 33658 30144 33934
rect 30196 33924 30248 33930
rect 30196 33866 30248 33872
rect 30104 33652 30156 33658
rect 30104 33594 30156 33600
rect 30116 33522 30144 33594
rect 30208 33522 30236 33866
rect 30564 33856 30616 33862
rect 30564 33798 30616 33804
rect 30380 33584 30432 33590
rect 30380 33526 30432 33532
rect 30104 33516 30156 33522
rect 30104 33458 30156 33464
rect 30196 33516 30248 33522
rect 30196 33458 30248 33464
rect 29184 33108 29236 33114
rect 29184 33050 29236 33056
rect 29736 32972 29788 32978
rect 29736 32914 29788 32920
rect 29092 32428 29144 32434
rect 29092 32370 29144 32376
rect 29748 31822 29776 32914
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 28908 31680 28960 31686
rect 28908 31622 28960 31628
rect 28724 30660 28776 30666
rect 28724 30602 28776 30608
rect 28736 30394 28764 30602
rect 28816 30592 28868 30598
rect 28816 30534 28868 30540
rect 28724 30388 28776 30394
rect 28724 30330 28776 30336
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28632 29776 28684 29782
rect 28632 29718 28684 29724
rect 28736 29714 28764 29990
rect 28724 29708 28776 29714
rect 28724 29650 28776 29656
rect 28632 29640 28684 29646
rect 28632 29582 28684 29588
rect 28644 29306 28672 29582
rect 28632 29300 28684 29306
rect 28632 29242 28684 29248
rect 28540 29232 28592 29238
rect 28368 29180 28540 29186
rect 28368 29174 28592 29180
rect 28264 29164 28316 29170
rect 28264 29106 28316 29112
rect 28368 29158 28580 29174
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28276 28082 28304 28494
rect 28368 28150 28396 29158
rect 28448 29096 28500 29102
rect 28448 29038 28500 29044
rect 28540 29096 28592 29102
rect 28540 29038 28592 29044
rect 28356 28144 28408 28150
rect 28356 28086 28408 28092
rect 28460 28082 28488 29038
rect 28264 28076 28316 28082
rect 28264 28018 28316 28024
rect 28448 28076 28500 28082
rect 28448 28018 28500 28024
rect 28552 27606 28580 29038
rect 28828 28558 28856 30534
rect 28920 30326 28948 31622
rect 29748 31498 29776 31758
rect 30104 31680 30156 31686
rect 30104 31622 30156 31628
rect 29656 31470 29776 31498
rect 29368 30864 29420 30870
rect 29368 30806 29420 30812
rect 29184 30728 29236 30734
rect 29184 30670 29236 30676
rect 29000 30660 29052 30666
rect 29052 30620 29132 30648
rect 29000 30602 29052 30608
rect 28908 30320 28960 30326
rect 28908 30262 28960 30268
rect 28920 29714 28948 30262
rect 28908 29708 28960 29714
rect 28908 29650 28960 29656
rect 28908 29504 28960 29510
rect 28908 29446 28960 29452
rect 28816 28552 28868 28558
rect 28816 28494 28868 28500
rect 28540 27600 28592 27606
rect 28540 27542 28592 27548
rect 27712 27464 27764 27470
rect 27712 27406 27764 27412
rect 27896 27464 27948 27470
rect 27896 27406 27948 27412
rect 28172 27464 28224 27470
rect 28224 27424 28304 27452
rect 28172 27406 28224 27412
rect 27620 26920 27672 26926
rect 27620 26862 27672 26868
rect 26424 26784 26476 26790
rect 26424 26726 26476 26732
rect 26516 26784 26568 26790
rect 26516 26726 26568 26732
rect 26240 26376 26292 26382
rect 26292 26336 26464 26364
rect 26240 26318 26292 26324
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 26332 25832 26384 25838
rect 26332 25774 26384 25780
rect 26344 25430 26372 25774
rect 26332 25424 26384 25430
rect 26332 25366 26384 25372
rect 26240 25356 26292 25362
rect 26240 25298 26292 25304
rect 25872 25288 25924 25294
rect 25872 25230 25924 25236
rect 25884 24614 25912 25230
rect 26252 24834 26280 25298
rect 25976 24818 26280 24834
rect 25964 24812 26280 24818
rect 26016 24806 26280 24812
rect 25964 24754 26016 24760
rect 25412 24608 25464 24614
rect 25412 24550 25464 24556
rect 25872 24608 25924 24614
rect 25872 24550 25924 24556
rect 25424 24206 25452 24550
rect 26252 24410 26280 24806
rect 26344 24750 26372 25366
rect 26436 24818 26464 26336
rect 26528 25974 26556 26726
rect 27724 26586 27752 27406
rect 27908 27062 27936 27406
rect 28172 27328 28224 27334
rect 28172 27270 28224 27276
rect 27896 27056 27948 27062
rect 27896 26998 27948 27004
rect 27908 26586 27936 26998
rect 28184 26994 28212 27270
rect 28276 26994 28304 27424
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 28264 26988 28316 26994
rect 28264 26930 28316 26936
rect 27712 26580 27764 26586
rect 27712 26522 27764 26528
rect 27896 26580 27948 26586
rect 27896 26522 27948 26528
rect 27160 26376 27212 26382
rect 27160 26318 27212 26324
rect 28540 26376 28592 26382
rect 28540 26318 28592 26324
rect 26516 25968 26568 25974
rect 26516 25910 26568 25916
rect 26528 25294 26556 25910
rect 27172 25498 27200 26318
rect 27160 25492 27212 25498
rect 27160 25434 27212 25440
rect 26516 25288 26568 25294
rect 26516 25230 26568 25236
rect 27804 25288 27856 25294
rect 27804 25230 27856 25236
rect 27620 25220 27672 25226
rect 27620 25162 27672 25168
rect 26516 25152 26568 25158
rect 26516 25094 26568 25100
rect 26528 24886 26556 25094
rect 27632 24954 27660 25162
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 26516 24880 26568 24886
rect 26516 24822 26568 24828
rect 26424 24812 26476 24818
rect 26424 24754 26476 24760
rect 26332 24744 26384 24750
rect 26332 24686 26384 24692
rect 26240 24404 26292 24410
rect 26240 24346 26292 24352
rect 26344 24274 26372 24686
rect 26528 24410 26556 24822
rect 26516 24404 26568 24410
rect 26516 24346 26568 24352
rect 26332 24268 26384 24274
rect 26332 24210 26384 24216
rect 27632 24206 27660 24890
rect 27816 24410 27844 25230
rect 27896 25152 27948 25158
rect 27896 25094 27948 25100
rect 27908 24818 27936 25094
rect 28552 24954 28580 26318
rect 28816 25900 28868 25906
rect 28816 25842 28868 25848
rect 28828 25226 28856 25842
rect 28816 25220 28868 25226
rect 28816 25162 28868 25168
rect 28540 24948 28592 24954
rect 28540 24890 28592 24896
rect 27896 24812 27948 24818
rect 27896 24754 27948 24760
rect 28540 24812 28592 24818
rect 28540 24754 28592 24760
rect 28552 24410 28580 24754
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 28540 24404 28592 24410
rect 28540 24346 28592 24352
rect 25412 24200 25464 24206
rect 25412 24142 25464 24148
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 28724 24200 28776 24206
rect 28920 24177 28948 29446
rect 29104 27334 29132 30620
rect 29196 30394 29224 30670
rect 29184 30388 29236 30394
rect 29184 30330 29236 30336
rect 29380 30258 29408 30806
rect 29656 30734 29684 31470
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 29748 30938 29776 31282
rect 30116 30938 30144 31622
rect 30208 31482 30236 33458
rect 30392 32842 30420 33526
rect 30576 33522 30604 33798
rect 30564 33516 30616 33522
rect 30564 33458 30616 33464
rect 30576 33318 30604 33458
rect 30564 33312 30616 33318
rect 30564 33254 30616 33260
rect 30576 33114 30604 33254
rect 30564 33108 30616 33114
rect 30564 33050 30616 33056
rect 30380 32836 30432 32842
rect 30380 32778 30432 32784
rect 30564 32836 30616 32842
rect 30564 32778 30616 32784
rect 30392 32570 30420 32778
rect 30380 32564 30432 32570
rect 30380 32506 30432 32512
rect 30576 32434 30604 32778
rect 30840 32768 30892 32774
rect 30840 32710 30892 32716
rect 30852 32434 30880 32710
rect 31036 32570 31064 33934
rect 31220 32910 31248 34070
rect 31668 33992 31720 33998
rect 31668 33934 31720 33940
rect 31392 33312 31444 33318
rect 31392 33254 31444 33260
rect 31404 33114 31432 33254
rect 31392 33108 31444 33114
rect 31392 33050 31444 33056
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31024 32564 31076 32570
rect 31024 32506 31076 32512
rect 30564 32428 30616 32434
rect 30564 32370 30616 32376
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 30944 32298 30972 32370
rect 31680 32366 31708 33934
rect 31668 32360 31720 32366
rect 31668 32302 31720 32308
rect 30932 32292 30984 32298
rect 30932 32234 30984 32240
rect 30748 32224 30800 32230
rect 30748 32166 30800 32172
rect 31680 32178 31708 32302
rect 30760 31822 30788 32166
rect 31680 32150 31800 32178
rect 31772 32026 31800 32150
rect 31668 32020 31720 32026
rect 31668 31962 31720 31968
rect 31760 32020 31812 32026
rect 31760 31962 31812 31968
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30288 31748 30340 31754
rect 30288 31690 30340 31696
rect 30196 31476 30248 31482
rect 30196 31418 30248 31424
rect 29736 30932 29788 30938
rect 29736 30874 29788 30880
rect 30104 30932 30156 30938
rect 30104 30874 30156 30880
rect 30208 30734 30236 31418
rect 30300 31414 30328 31690
rect 30288 31408 30340 31414
rect 30288 31350 30340 31356
rect 30300 30734 30328 31350
rect 31680 31346 31708 31962
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 31300 31136 31352 31142
rect 31300 31078 31352 31084
rect 29644 30728 29696 30734
rect 29644 30670 29696 30676
rect 30196 30728 30248 30734
rect 30196 30670 30248 30676
rect 30288 30728 30340 30734
rect 30288 30670 30340 30676
rect 29368 30252 29420 30258
rect 29368 30194 29420 30200
rect 29380 29170 29408 30194
rect 29460 30184 29512 30190
rect 29460 30126 29512 30132
rect 29472 29850 29500 30126
rect 30012 30116 30064 30122
rect 30012 30058 30064 30064
rect 29460 29844 29512 29850
rect 29460 29786 29512 29792
rect 29472 29238 29500 29786
rect 29644 29504 29696 29510
rect 29644 29446 29696 29452
rect 29460 29232 29512 29238
rect 29460 29174 29512 29180
rect 29656 29170 29684 29446
rect 29368 29164 29420 29170
rect 29368 29106 29420 29112
rect 29644 29164 29696 29170
rect 29644 29106 29696 29112
rect 29276 28688 29328 28694
rect 29276 28630 29328 28636
rect 29288 27946 29316 28630
rect 30024 28082 30052 30058
rect 30300 29238 30328 30670
rect 31312 30666 31340 31078
rect 31300 30660 31352 30666
rect 31300 30602 31352 30608
rect 31392 30660 31444 30666
rect 31392 30602 31444 30608
rect 30564 29776 30616 29782
rect 30564 29718 30616 29724
rect 30288 29232 30340 29238
rect 30288 29174 30340 29180
rect 30380 28416 30432 28422
rect 30380 28358 30432 28364
rect 30392 28082 30420 28358
rect 30012 28076 30064 28082
rect 30012 28018 30064 28024
rect 30196 28076 30248 28082
rect 30196 28018 30248 28024
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 29184 27940 29236 27946
rect 29184 27882 29236 27888
rect 29276 27940 29328 27946
rect 29276 27882 29328 27888
rect 29196 27470 29224 27882
rect 29552 27872 29604 27878
rect 29552 27814 29604 27820
rect 29184 27464 29236 27470
rect 29184 27406 29236 27412
rect 29092 27328 29144 27334
rect 29092 27270 29144 27276
rect 29460 27328 29512 27334
rect 29460 27270 29512 27276
rect 29000 26988 29052 26994
rect 29000 26930 29052 26936
rect 29012 26586 29040 26930
rect 29000 26580 29052 26586
rect 29000 26522 29052 26528
rect 29000 26376 29052 26382
rect 29000 26318 29052 26324
rect 29012 25498 29040 26318
rect 29368 25832 29420 25838
rect 29368 25774 29420 25780
rect 29184 25696 29236 25702
rect 29184 25638 29236 25644
rect 29000 25492 29052 25498
rect 29000 25434 29052 25440
rect 29000 25356 29052 25362
rect 29000 25298 29052 25304
rect 29012 24750 29040 25298
rect 29000 24744 29052 24750
rect 29000 24686 29052 24692
rect 28724 24142 28776 24148
rect 28906 24168 28962 24177
rect 28736 23866 28764 24142
rect 28906 24103 28962 24112
rect 28724 23860 28776 23866
rect 28724 23802 28776 23808
rect 25964 23724 26016 23730
rect 25964 23666 26016 23672
rect 26240 23724 26292 23730
rect 26976 23724 27028 23730
rect 26292 23684 26372 23712
rect 26240 23666 26292 23672
rect 25976 23050 26004 23666
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26252 23186 26280 23462
rect 26344 23186 26372 23684
rect 26976 23666 27028 23672
rect 26240 23180 26292 23186
rect 26240 23122 26292 23128
rect 26332 23180 26384 23186
rect 26332 23122 26384 23128
rect 25964 23044 26016 23050
rect 25964 22986 26016 22992
rect 25688 22976 25740 22982
rect 25688 22918 25740 22924
rect 25700 22778 25728 22918
rect 26344 22778 26372 23122
rect 26792 23112 26844 23118
rect 26988 23100 27016 23666
rect 26844 23072 27016 23100
rect 26792 23054 26844 23060
rect 25688 22772 25740 22778
rect 25688 22714 25740 22720
rect 26332 22772 26384 22778
rect 26332 22714 26384 22720
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 26516 22568 26568 22574
rect 26516 22510 26568 22516
rect 25792 22030 25820 22510
rect 26528 22098 26556 22510
rect 26988 22166 27016 23072
rect 27988 22636 28040 22642
rect 27988 22578 28040 22584
rect 27712 22568 27764 22574
rect 27712 22510 27764 22516
rect 26976 22160 27028 22166
rect 26976 22102 27028 22108
rect 26516 22092 26568 22098
rect 26516 22034 26568 22040
rect 25780 22024 25832 22030
rect 25780 21966 25832 21972
rect 26792 22024 26844 22030
rect 26792 21966 26844 21972
rect 25228 21956 25280 21962
rect 25228 21898 25280 21904
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25240 21350 25268 21898
rect 26240 21548 26292 21554
rect 26240 21490 26292 21496
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 25504 21344 25556 21350
rect 25504 21286 25556 21292
rect 25136 20800 25188 20806
rect 25136 20742 25188 20748
rect 25148 20398 25176 20742
rect 25136 20392 25188 20398
rect 25136 20334 25188 20340
rect 25148 19854 25176 20334
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25044 18624 25096 18630
rect 25044 18566 25096 18572
rect 25056 17660 25084 18566
rect 25148 18086 25176 19790
rect 25240 19786 25268 21286
rect 25516 20466 25544 21286
rect 25504 20460 25556 20466
rect 25504 20402 25556 20408
rect 26252 20058 26280 21490
rect 26700 21344 26752 21350
rect 26700 21286 26752 21292
rect 26712 20874 26740 21286
rect 26700 20868 26752 20874
rect 26700 20810 26752 20816
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25596 19916 25648 19922
rect 25596 19858 25648 19864
rect 25228 19780 25280 19786
rect 25228 19722 25280 19728
rect 25608 19514 25636 19858
rect 25596 19508 25648 19514
rect 25596 19450 25648 19456
rect 25596 18692 25648 18698
rect 25596 18634 25648 18640
rect 25608 18426 25636 18634
rect 25596 18420 25648 18426
rect 25596 18362 25648 18368
rect 25792 18290 25820 19926
rect 25964 19712 26016 19718
rect 25964 19654 26016 19660
rect 25976 18970 26004 19654
rect 26240 19372 26292 19378
rect 26240 19314 26292 19320
rect 25964 18964 26016 18970
rect 25964 18906 26016 18912
rect 25976 18290 26004 18906
rect 25780 18284 25832 18290
rect 25780 18226 25832 18232
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25136 18080 25188 18086
rect 25136 18022 25188 18028
rect 25872 18080 25924 18086
rect 25872 18022 25924 18028
rect 25504 17808 25556 17814
rect 25504 17750 25556 17756
rect 25136 17672 25188 17678
rect 25056 17632 25136 17660
rect 25136 17614 25188 17620
rect 25228 17604 25280 17610
rect 25412 17604 25464 17610
rect 25228 17546 25280 17552
rect 25332 17564 25412 17592
rect 25136 17332 25188 17338
rect 25136 17274 25188 17280
rect 24952 17128 25004 17134
rect 24952 17070 25004 17076
rect 24860 17060 24912 17066
rect 24860 17002 24912 17008
rect 23664 16652 23716 16658
rect 23664 16594 23716 16600
rect 24676 16652 24728 16658
rect 24676 16594 24728 16600
rect 23572 16108 23624 16114
rect 23572 16050 23624 16056
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 23112 15700 23164 15706
rect 23112 15642 23164 15648
rect 23480 15700 23532 15706
rect 23480 15642 23532 15648
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22652 15496 22704 15502
rect 22652 15438 22704 15444
rect 20812 14272 20864 14278
rect 20812 14214 20864 14220
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20628 13524 20680 13530
rect 20628 13466 20680 13472
rect 20732 13394 20760 13874
rect 20720 13388 20772 13394
rect 20720 13330 20772 13336
rect 19800 13320 19852 13326
rect 19800 13262 19852 13268
rect 20444 13320 20496 13326
rect 20444 13262 20496 13268
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 20732 12986 20760 13330
rect 20824 13326 20852 14214
rect 21192 13870 21220 15438
rect 21456 15428 21508 15434
rect 21456 15370 21508 15376
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21272 15020 21324 15026
rect 21272 14962 21324 14968
rect 21284 14618 21312 14962
rect 21272 14612 21324 14618
rect 21272 14554 21324 14560
rect 21376 14346 21404 15302
rect 21468 14822 21496 15370
rect 22112 15162 22140 15438
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22744 15156 22796 15162
rect 22744 15098 22796 15104
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14396 21496 14758
rect 22190 14512 22246 14521
rect 22190 14447 22246 14456
rect 21548 14408 21600 14414
rect 21468 14368 21548 14396
rect 21364 14340 21416 14346
rect 21364 14282 21416 14288
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21180 13864 21232 13870
rect 21180 13806 21232 13812
rect 21284 13530 21312 14214
rect 21376 14006 21404 14282
rect 21364 14000 21416 14006
rect 21364 13942 21416 13948
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21376 13326 21404 13942
rect 20812 13320 20864 13326
rect 20812 13262 20864 13268
rect 20904 13320 20956 13326
rect 20904 13262 20956 13268
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 20720 12980 20772 12986
rect 20720 12922 20772 12928
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20272 12442 20300 12786
rect 20536 12776 20588 12782
rect 20536 12718 20588 12724
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20260 12436 20312 12442
rect 20260 12378 20312 12384
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 20272 11762 20300 12378
rect 20456 12306 20484 12582
rect 20548 12442 20576 12718
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20444 12300 20496 12306
rect 20444 12242 20496 12248
rect 20260 11756 20312 11762
rect 20260 11698 20312 11704
rect 20548 11558 20576 12378
rect 20916 12374 20944 13262
rect 20904 12368 20956 12374
rect 20904 12310 20956 12316
rect 21468 12238 21496 14368
rect 21548 14350 21600 14356
rect 22204 13938 22232 14447
rect 22756 13938 22784 15098
rect 23584 15094 23612 16050
rect 23664 15496 23716 15502
rect 23664 15438 23716 15444
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 22928 15020 22980 15026
rect 22928 14962 22980 14968
rect 22940 14074 22968 14962
rect 23572 14408 23624 14414
rect 23676 14396 23704 15438
rect 24688 15094 24716 16594
rect 25148 16590 25176 17274
rect 24952 16584 25004 16590
rect 24952 16526 25004 16532
rect 25136 16584 25188 16590
rect 25136 16526 25188 16532
rect 24964 16250 24992 16526
rect 24952 16244 25004 16250
rect 24952 16186 25004 16192
rect 25148 16114 25176 16526
rect 25136 16108 25188 16114
rect 25136 16050 25188 16056
rect 25240 15434 25268 17546
rect 25332 17270 25360 17564
rect 25412 17546 25464 17552
rect 25320 17264 25372 17270
rect 25320 17206 25372 17212
rect 25332 16590 25360 17206
rect 25516 16590 25544 17750
rect 25884 17610 25912 18022
rect 25976 17882 26004 18226
rect 25964 17876 26016 17882
rect 25964 17818 26016 17824
rect 25872 17604 25924 17610
rect 25872 17546 25924 17552
rect 25596 16992 25648 16998
rect 25596 16934 25648 16940
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25504 16584 25556 16590
rect 25504 16526 25556 16532
rect 25332 15978 25360 16526
rect 25412 16516 25464 16522
rect 25412 16458 25464 16464
rect 25424 15978 25452 16458
rect 25320 15972 25372 15978
rect 25320 15914 25372 15920
rect 25412 15972 25464 15978
rect 25412 15914 25464 15920
rect 25320 15496 25372 15502
rect 25320 15438 25372 15444
rect 25228 15428 25280 15434
rect 25228 15370 25280 15376
rect 25332 15162 25360 15438
rect 25516 15162 25544 16526
rect 25608 16182 25636 16934
rect 25596 16176 25648 16182
rect 25596 16118 25648 16124
rect 25884 16114 25912 17546
rect 25976 17338 26004 17818
rect 26148 17536 26200 17542
rect 26148 17478 26200 17484
rect 25964 17332 26016 17338
rect 25964 17274 26016 17280
rect 26160 17202 26188 17478
rect 26148 17196 26200 17202
rect 26148 17138 26200 17144
rect 25872 16108 25924 16114
rect 25872 16050 25924 16056
rect 26252 15910 26280 19314
rect 26804 17678 26832 21966
rect 27344 21548 27396 21554
rect 27344 21490 27396 21496
rect 27356 19854 27384 21490
rect 27528 21480 27580 21486
rect 27528 21422 27580 21428
rect 27540 20874 27568 21422
rect 27724 20942 27752 22510
rect 28000 21690 28028 22578
rect 28540 22024 28592 22030
rect 28540 21966 28592 21972
rect 28552 21690 28580 21966
rect 27988 21684 28040 21690
rect 27988 21626 28040 21632
rect 28540 21684 28592 21690
rect 28540 21626 28592 21632
rect 28816 21548 28868 21554
rect 28816 21490 28868 21496
rect 28172 21480 28224 21486
rect 28172 21422 28224 21428
rect 28448 21480 28500 21486
rect 28448 21422 28500 21428
rect 28632 21480 28684 21486
rect 28632 21422 28684 21428
rect 28080 21412 28132 21418
rect 28080 21354 28132 21360
rect 27712 20936 27764 20942
rect 27712 20878 27764 20884
rect 27528 20868 27580 20874
rect 27528 20810 27580 20816
rect 27540 20466 27568 20810
rect 27724 20534 27752 20878
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 27712 20528 27764 20534
rect 27712 20470 27764 20476
rect 27528 20460 27580 20466
rect 27528 20402 27580 20408
rect 27724 20398 27752 20470
rect 28000 20466 28028 20742
rect 27988 20460 28040 20466
rect 27988 20402 28040 20408
rect 27712 20392 27764 20398
rect 27712 20334 27764 20340
rect 27344 19848 27396 19854
rect 27344 19790 27396 19796
rect 27160 19780 27212 19786
rect 27160 19722 27212 19728
rect 26792 17672 26844 17678
rect 26792 17614 26844 17620
rect 26516 17604 26568 17610
rect 26516 17546 26568 17552
rect 26528 17202 26556 17546
rect 27172 17270 27200 19722
rect 27344 19372 27396 19378
rect 27724 19360 27752 20334
rect 28000 19922 28028 20402
rect 27988 19916 28040 19922
rect 27988 19858 28040 19864
rect 28092 19802 28120 21354
rect 28184 21146 28212 21422
rect 28172 21140 28224 21146
rect 28172 21082 28224 21088
rect 28356 21072 28408 21078
rect 28356 21014 28408 21020
rect 28368 20058 28396 21014
rect 28460 20262 28488 21422
rect 28644 21078 28672 21422
rect 28632 21072 28684 21078
rect 28632 21014 28684 21020
rect 28644 20942 28672 21014
rect 28632 20936 28684 20942
rect 28632 20878 28684 20884
rect 28540 20800 28592 20806
rect 28540 20742 28592 20748
rect 28552 20262 28580 20742
rect 28632 20324 28684 20330
rect 28632 20266 28684 20272
rect 28448 20256 28500 20262
rect 28448 20198 28500 20204
rect 28540 20256 28592 20262
rect 28540 20198 28592 20204
rect 28356 20052 28408 20058
rect 28356 19994 28408 20000
rect 28552 19854 28580 20198
rect 28644 20058 28672 20266
rect 28632 20052 28684 20058
rect 28632 19994 28684 20000
rect 27344 19314 27396 19320
rect 27540 19332 27752 19360
rect 28000 19774 28120 19802
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28540 19848 28592 19854
rect 28540 19790 28592 19796
rect 27252 19168 27304 19174
rect 27252 19110 27304 19116
rect 27264 18290 27292 19110
rect 27252 18284 27304 18290
rect 27252 18226 27304 18232
rect 27356 17882 27384 19314
rect 27540 18766 27568 19332
rect 27528 18760 27580 18766
rect 27528 18702 27580 18708
rect 27540 18358 27568 18702
rect 27712 18624 27764 18630
rect 27712 18566 27764 18572
rect 27528 18352 27580 18358
rect 27528 18294 27580 18300
rect 27344 17876 27396 17882
rect 27344 17818 27396 17824
rect 27724 17610 27752 18566
rect 27712 17604 27764 17610
rect 27712 17546 27764 17552
rect 27160 17264 27212 17270
rect 27160 17206 27212 17212
rect 27528 17264 27580 17270
rect 27528 17206 27580 17212
rect 26516 17196 26568 17202
rect 26516 17138 26568 17144
rect 27252 17196 27304 17202
rect 27252 17138 27304 17144
rect 27160 16516 27212 16522
rect 27160 16458 27212 16464
rect 27172 16250 27200 16458
rect 27160 16244 27212 16250
rect 27160 16186 27212 16192
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 27264 15570 27292 17138
rect 27344 16992 27396 16998
rect 27344 16934 27396 16940
rect 27356 16114 27384 16934
rect 27540 16454 27568 17206
rect 27528 16448 27580 16454
rect 27528 16390 27580 16396
rect 27540 16114 27568 16390
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27528 16108 27580 16114
rect 27528 16050 27580 16056
rect 27252 15564 27304 15570
rect 27252 15506 27304 15512
rect 25872 15428 25924 15434
rect 25872 15370 25924 15376
rect 25320 15156 25372 15162
rect 25320 15098 25372 15104
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25884 15094 25912 15370
rect 24676 15088 24728 15094
rect 24676 15030 24728 15036
rect 25872 15088 25924 15094
rect 25872 15030 25924 15036
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24044 14618 24072 14962
rect 24032 14612 24084 14618
rect 24032 14554 24084 14560
rect 24688 14482 24716 15030
rect 26332 15020 26384 15026
rect 26332 14962 26384 14968
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 24124 14476 24176 14482
rect 24124 14418 24176 14424
rect 24676 14476 24728 14482
rect 24676 14418 24728 14424
rect 23624 14368 23704 14396
rect 23572 14350 23624 14356
rect 22928 14068 22980 14074
rect 22928 14010 22980 14016
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22376 13932 22428 13938
rect 22376 13874 22428 13880
rect 22744 13932 22796 13938
rect 22744 13874 22796 13880
rect 22008 13864 22060 13870
rect 22060 13812 22140 13818
rect 22008 13806 22140 13812
rect 22020 13790 22140 13806
rect 22112 13394 22140 13790
rect 22100 13388 22152 13394
rect 22100 13330 22152 13336
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22296 12850 22324 13194
rect 22388 12986 22416 13874
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22480 13530 22508 13806
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22468 13320 22520 13326
rect 22468 13262 22520 13268
rect 22376 12980 22428 12986
rect 22376 12922 22428 12928
rect 22480 12850 22508 13262
rect 22756 12850 22784 13874
rect 23676 13190 23704 14368
rect 23940 14340 23992 14346
rect 23940 14282 23992 14288
rect 23952 14006 23980 14282
rect 24136 14074 24164 14418
rect 25780 14408 25832 14414
rect 25780 14350 25832 14356
rect 25228 14340 25280 14346
rect 25228 14282 25280 14288
rect 25240 14074 25268 14282
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 25228 14068 25280 14074
rect 25228 14010 25280 14016
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 25792 13938 25820 14350
rect 26344 14278 26372 14962
rect 26332 14272 26384 14278
rect 26332 14214 26384 14220
rect 23756 13932 23808 13938
rect 23756 13874 23808 13880
rect 25596 13932 25648 13938
rect 25596 13874 25648 13880
rect 25780 13932 25832 13938
rect 25780 13874 25832 13880
rect 23664 13184 23716 13190
rect 23664 13126 23716 13132
rect 23676 12850 23704 13126
rect 23768 12986 23796 13874
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 23848 13728 23900 13734
rect 23848 13670 23900 13676
rect 23860 13326 23888 13670
rect 23848 13320 23900 13326
rect 23848 13262 23900 13268
rect 23940 13320 23992 13326
rect 23940 13262 23992 13268
rect 23756 12980 23808 12986
rect 23756 12922 23808 12928
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 22744 12844 22796 12850
rect 22744 12786 22796 12792
rect 23664 12844 23716 12850
rect 23664 12786 23716 12792
rect 22100 12708 22152 12714
rect 22100 12650 22152 12656
rect 22112 12306 22140 12650
rect 22480 12374 22508 12786
rect 22468 12368 22520 12374
rect 22468 12310 22520 12316
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 22756 12238 22784 12786
rect 23388 12776 23440 12782
rect 23388 12718 23440 12724
rect 20812 12232 20864 12238
rect 20812 12174 20864 12180
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 22744 12232 22796 12238
rect 22744 12174 22796 12180
rect 23296 12232 23348 12238
rect 23400 12220 23428 12718
rect 23480 12640 23532 12646
rect 23480 12582 23532 12588
rect 23492 12238 23520 12582
rect 23348 12192 23428 12220
rect 23480 12232 23532 12238
rect 23296 12174 23348 12180
rect 23480 12174 23532 12180
rect 20824 11898 20852 12174
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 23676 11762 23704 12786
rect 23952 12714 23980 13262
rect 24676 13252 24728 13258
rect 24676 13194 24728 13200
rect 24688 12986 24716 13194
rect 24872 13190 24900 13806
rect 25608 13530 25636 13874
rect 26344 13870 26372 14214
rect 26436 14006 26464 14962
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26332 13864 26384 13870
rect 26332 13806 26384 13812
rect 25596 13524 25648 13530
rect 25596 13466 25648 13472
rect 25964 13320 26016 13326
rect 26016 13280 26280 13308
rect 25964 13262 26016 13268
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24676 12980 24728 12986
rect 24676 12922 24728 12928
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 23940 12708 23992 12714
rect 23940 12650 23992 12656
rect 23664 11756 23716 11762
rect 23664 11698 23716 11704
rect 23952 11694 23980 12650
rect 24044 12374 24072 12786
rect 24780 12442 24808 12786
rect 26252 12714 26280 13280
rect 26344 12850 26372 13806
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26436 12730 26464 13942
rect 26700 13320 26752 13326
rect 26700 13262 26752 13268
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26344 12714 26556 12730
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26332 12708 26556 12714
rect 26384 12702 26556 12708
rect 26332 12650 26384 12656
rect 24768 12436 24820 12442
rect 24768 12378 24820 12384
rect 26252 12374 26280 12650
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 24032 12368 24084 12374
rect 24032 12310 24084 12316
rect 26240 12368 26292 12374
rect 26240 12310 26292 12316
rect 24044 11898 24072 12310
rect 26436 12238 26464 12582
rect 26528 12374 26556 12702
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26712 12170 26740 13262
rect 26804 12306 26832 13262
rect 27264 13190 27292 15506
rect 27540 15434 27568 16050
rect 27896 15904 27948 15910
rect 27896 15846 27948 15852
rect 27804 15700 27856 15706
rect 27804 15642 27856 15648
rect 27712 15496 27764 15502
rect 27712 15438 27764 15444
rect 27528 15428 27580 15434
rect 27528 15370 27580 15376
rect 27540 15094 27568 15370
rect 27620 15360 27672 15366
rect 27620 15302 27672 15308
rect 27528 15088 27580 15094
rect 27528 15030 27580 15036
rect 27344 14816 27396 14822
rect 27344 14758 27396 14764
rect 27356 13462 27384 14758
rect 27540 14346 27568 15030
rect 27632 15026 27660 15302
rect 27724 15162 27752 15438
rect 27712 15156 27764 15162
rect 27712 15098 27764 15104
rect 27620 15020 27672 15026
rect 27620 14962 27672 14968
rect 27632 14618 27660 14962
rect 27620 14612 27672 14618
rect 27620 14554 27672 14560
rect 27724 14346 27752 15098
rect 27816 14618 27844 15642
rect 27908 15570 27936 15846
rect 27896 15564 27948 15570
rect 27896 15506 27948 15512
rect 27804 14612 27856 14618
rect 27804 14554 27856 14560
rect 27908 14346 27936 15506
rect 28000 14521 28028 19774
rect 28276 19514 28304 19790
rect 28264 19508 28316 19514
rect 28264 19450 28316 19456
rect 28172 19372 28224 19378
rect 28172 19314 28224 19320
rect 28264 19372 28316 19378
rect 28264 19314 28316 19320
rect 28080 18692 28132 18698
rect 28080 18634 28132 18640
rect 28092 17882 28120 18634
rect 28184 18630 28212 19314
rect 28276 18766 28304 19314
rect 28356 19304 28408 19310
rect 28356 19246 28408 19252
rect 28368 18766 28396 19246
rect 28724 19168 28776 19174
rect 28724 19110 28776 19116
rect 28264 18760 28316 18766
rect 28264 18702 28316 18708
rect 28356 18760 28408 18766
rect 28356 18702 28408 18708
rect 28172 18624 28224 18630
rect 28172 18566 28224 18572
rect 28080 17876 28132 17882
rect 28080 17818 28132 17824
rect 28276 17814 28304 18702
rect 28368 18426 28396 18702
rect 28736 18698 28764 19110
rect 28828 18970 28856 21490
rect 28920 21418 28948 24103
rect 29012 23644 29040 24686
rect 29196 24410 29224 25638
rect 29380 25498 29408 25774
rect 29276 25492 29328 25498
rect 29276 25434 29328 25440
rect 29368 25492 29420 25498
rect 29368 25434 29420 25440
rect 29288 24614 29316 25434
rect 29368 25220 29420 25226
rect 29368 25162 29420 25168
rect 29276 24608 29328 24614
rect 29276 24550 29328 24556
rect 29184 24404 29236 24410
rect 29184 24346 29236 24352
rect 29196 23866 29224 24346
rect 29288 24206 29316 24550
rect 29380 24342 29408 25162
rect 29368 24336 29420 24342
rect 29368 24278 29420 24284
rect 29276 24200 29328 24206
rect 29276 24142 29328 24148
rect 29184 23860 29236 23866
rect 29184 23802 29236 23808
rect 29472 23730 29500 27270
rect 29564 26994 29592 27814
rect 30024 27606 30052 28018
rect 30012 27600 30064 27606
rect 30012 27542 30064 27548
rect 30208 27538 30236 28018
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30484 27606 30512 27950
rect 30472 27600 30524 27606
rect 30472 27542 30524 27548
rect 29644 27532 29696 27538
rect 29644 27474 29696 27480
rect 30196 27532 30248 27538
rect 30196 27474 30248 27480
rect 29552 26988 29604 26994
rect 29552 26930 29604 26936
rect 29460 23724 29512 23730
rect 29460 23666 29512 23672
rect 29092 23656 29144 23662
rect 29012 23616 29092 23644
rect 29012 23118 29040 23616
rect 29092 23598 29144 23604
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29092 23044 29144 23050
rect 29092 22986 29144 22992
rect 29104 22234 29132 22986
rect 29092 22228 29144 22234
rect 29092 22170 29144 22176
rect 29000 22024 29052 22030
rect 29000 21966 29052 21972
rect 28908 21412 28960 21418
rect 28908 21354 28960 21360
rect 29012 20534 29040 21966
rect 29104 20602 29132 22170
rect 29564 22094 29592 26930
rect 29656 26042 29684 27474
rect 29736 27464 29788 27470
rect 29736 27406 29788 27412
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 29748 27130 29776 27406
rect 29736 27124 29788 27130
rect 29736 27066 29788 27072
rect 29932 27062 29960 27406
rect 29920 27056 29972 27062
rect 29920 26998 29972 27004
rect 30024 26994 30052 27406
rect 30196 27328 30248 27334
rect 30196 27270 30248 27276
rect 30208 26994 30236 27270
rect 30288 27124 30340 27130
rect 30288 27066 30340 27072
rect 30380 27124 30432 27130
rect 30380 27066 30432 27072
rect 30012 26988 30064 26994
rect 30012 26930 30064 26936
rect 30196 26988 30248 26994
rect 30196 26930 30248 26936
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30116 26382 30144 26726
rect 30300 26382 30328 27066
rect 30392 26450 30420 27066
rect 30380 26444 30432 26450
rect 30380 26386 30432 26392
rect 30104 26376 30156 26382
rect 30104 26318 30156 26324
rect 30288 26376 30340 26382
rect 30288 26318 30340 26324
rect 30196 26308 30248 26314
rect 30196 26250 30248 26256
rect 29644 26036 29696 26042
rect 29644 25978 29696 25984
rect 30208 25974 30236 26250
rect 30196 25968 30248 25974
rect 30196 25910 30248 25916
rect 29828 25832 29880 25838
rect 29828 25774 29880 25780
rect 29840 25362 29868 25774
rect 29828 25356 29880 25362
rect 29828 25298 29880 25304
rect 30012 25152 30064 25158
rect 30012 25094 30064 25100
rect 30024 24750 30052 25094
rect 30300 24750 30328 26318
rect 30012 24744 30064 24750
rect 30012 24686 30064 24692
rect 30288 24744 30340 24750
rect 30288 24686 30340 24692
rect 30576 22778 30604 29718
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 30944 29306 30972 29582
rect 30932 29300 30984 29306
rect 30932 29242 30984 29248
rect 30748 28620 30800 28626
rect 30748 28562 30800 28568
rect 30656 28416 30708 28422
rect 30656 28358 30708 28364
rect 30668 28218 30696 28358
rect 30760 28218 30788 28562
rect 30656 28212 30708 28218
rect 30656 28154 30708 28160
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30944 28150 30972 29242
rect 31404 28558 31432 30602
rect 31852 30592 31904 30598
rect 31852 30534 31904 30540
rect 31864 29646 31892 30534
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 32220 29640 32272 29646
rect 32220 29582 32272 29588
rect 31760 29504 31812 29510
rect 31760 29446 31812 29452
rect 31772 29170 31800 29446
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 31668 28960 31720 28966
rect 31668 28902 31720 28908
rect 31680 28558 31708 28902
rect 31024 28552 31076 28558
rect 31024 28494 31076 28500
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31668 28552 31720 28558
rect 31668 28494 31720 28500
rect 30932 28144 30984 28150
rect 30932 28086 30984 28092
rect 30944 27878 30972 28086
rect 31036 28082 31064 28494
rect 32232 28490 32260 29582
rect 32324 28762 32352 35866
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34520 33448 34572 33454
rect 34520 33390 34572 33396
rect 34152 33380 34204 33386
rect 34152 33322 34204 33328
rect 33968 33312 34020 33318
rect 33968 33254 34020 33260
rect 33980 33114 34008 33254
rect 33968 33108 34020 33114
rect 33968 33050 34020 33056
rect 33692 32904 33744 32910
rect 33692 32846 33744 32852
rect 33784 32904 33836 32910
rect 33784 32846 33836 32852
rect 33704 32298 33732 32846
rect 33796 32570 33824 32846
rect 33784 32564 33836 32570
rect 33784 32506 33836 32512
rect 33876 32428 33928 32434
rect 33980 32416 34008 33050
rect 34060 32972 34112 32978
rect 34060 32914 34112 32920
rect 34072 32434 34100 32914
rect 34164 32842 34192 33322
rect 34532 33046 34560 33390
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34520 33040 34572 33046
rect 34520 32982 34572 32988
rect 34152 32836 34204 32842
rect 34152 32778 34204 32784
rect 33928 32388 34008 32416
rect 34060 32428 34112 32434
rect 33876 32370 33928 32376
rect 34060 32370 34112 32376
rect 34164 32314 34192 32778
rect 33692 32292 33744 32298
rect 33692 32234 33744 32240
rect 34072 32286 34192 32314
rect 34428 32360 34480 32366
rect 34428 32302 34480 32308
rect 32496 31816 32548 31822
rect 32496 31758 32548 31764
rect 32404 31748 32456 31754
rect 32404 31690 32456 31696
rect 32416 31482 32444 31690
rect 32404 31476 32456 31482
rect 32404 31418 32456 31424
rect 32508 30734 32536 31758
rect 33232 31340 33284 31346
rect 33232 31282 33284 31288
rect 33244 30938 33272 31282
rect 33232 30932 33284 30938
rect 33232 30874 33284 30880
rect 32496 30728 32548 30734
rect 32496 30670 32548 30676
rect 32772 29572 32824 29578
rect 32772 29514 32824 29520
rect 32784 29170 32812 29514
rect 33244 29170 33272 30874
rect 33968 30660 34020 30666
rect 33968 30602 34020 30608
rect 33980 30394 34008 30602
rect 34072 30598 34100 32286
rect 34440 32026 34468 32302
rect 34428 32020 34480 32026
rect 34428 31962 34480 31968
rect 34532 31634 34560 32982
rect 37648 32428 37700 32434
rect 37648 32370 37700 32376
rect 36268 32360 36320 32366
rect 36268 32302 36320 32308
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 36280 32026 36308 32302
rect 37188 32224 37240 32230
rect 37188 32166 37240 32172
rect 36268 32020 36320 32026
rect 36268 31962 36320 31968
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 35532 31816 35584 31822
rect 35532 31758 35584 31764
rect 36912 31816 36964 31822
rect 36912 31758 36964 31764
rect 34440 31606 34560 31634
rect 34440 31278 34468 31606
rect 34428 31272 34480 31278
rect 34428 31214 34480 31220
rect 34060 30592 34112 30598
rect 34060 30534 34112 30540
rect 33968 30388 34020 30394
rect 33968 30330 34020 30336
rect 33692 30320 33744 30326
rect 33692 30262 33744 30268
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 32864 29164 32916 29170
rect 32864 29106 32916 29112
rect 33232 29164 33284 29170
rect 33284 29124 33548 29152
rect 33232 29106 33284 29112
rect 32784 28762 32812 29106
rect 32312 28756 32364 28762
rect 32312 28698 32364 28704
rect 32772 28756 32824 28762
rect 32772 28698 32824 28704
rect 31300 28484 31352 28490
rect 31300 28426 31352 28432
rect 32036 28484 32088 28490
rect 32036 28426 32088 28432
rect 32220 28484 32272 28490
rect 32220 28426 32272 28432
rect 31024 28076 31076 28082
rect 31024 28018 31076 28024
rect 30932 27872 30984 27878
rect 30932 27814 30984 27820
rect 31036 27130 31064 28018
rect 31312 27334 31340 28426
rect 32048 28014 32076 28426
rect 32036 28008 32088 28014
rect 32036 27950 32088 27956
rect 32048 27470 32076 27950
rect 32232 27946 32260 28426
rect 32220 27940 32272 27946
rect 32220 27882 32272 27888
rect 32036 27464 32088 27470
rect 32036 27406 32088 27412
rect 31300 27328 31352 27334
rect 31300 27270 31352 27276
rect 31024 27124 31076 27130
rect 31024 27066 31076 27072
rect 31036 25770 31064 27066
rect 31312 27062 31340 27270
rect 31300 27056 31352 27062
rect 31300 26998 31352 27004
rect 31208 26308 31260 26314
rect 31208 26250 31260 26256
rect 31024 25764 31076 25770
rect 31024 25706 31076 25712
rect 30748 25696 30800 25702
rect 30748 25638 30800 25644
rect 30760 24818 30788 25638
rect 30840 25220 30892 25226
rect 30840 25162 30892 25168
rect 30748 24812 30800 24818
rect 30748 24754 30800 24760
rect 30852 24682 30880 25162
rect 30840 24676 30892 24682
rect 30840 24618 30892 24624
rect 31220 23322 31248 26250
rect 32048 26246 32076 27406
rect 32232 27130 32260 27882
rect 32588 27328 32640 27334
rect 32588 27270 32640 27276
rect 32220 27124 32272 27130
rect 32220 27066 32272 27072
rect 32600 26450 32628 27270
rect 32772 27124 32824 27130
rect 32772 27066 32824 27072
rect 32588 26444 32640 26450
rect 32588 26386 32640 26392
rect 32036 26240 32088 26246
rect 32036 26182 32088 26188
rect 31392 25900 31444 25906
rect 31392 25842 31444 25848
rect 31404 25498 31432 25842
rect 31392 25492 31444 25498
rect 31392 25434 31444 25440
rect 31944 24744 31996 24750
rect 31944 24686 31996 24692
rect 31760 24268 31812 24274
rect 31760 24210 31812 24216
rect 31772 24070 31800 24210
rect 31392 24064 31444 24070
rect 31392 24006 31444 24012
rect 31760 24064 31812 24070
rect 31760 24006 31812 24012
rect 31404 23798 31432 24006
rect 31392 23792 31444 23798
rect 31392 23734 31444 23740
rect 31208 23316 31260 23322
rect 31208 23258 31260 23264
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30576 22658 30604 22714
rect 30288 22636 30340 22642
rect 30288 22578 30340 22584
rect 30392 22630 30604 22658
rect 31116 22704 31168 22710
rect 31116 22646 31168 22652
rect 29564 22066 29684 22094
rect 29092 20596 29144 20602
rect 29092 20538 29144 20544
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29460 19712 29512 19718
rect 29460 19654 29512 19660
rect 29472 19378 29500 19654
rect 29656 19378 29684 22066
rect 30012 22024 30064 22030
rect 30012 21966 30064 21972
rect 29920 21548 29972 21554
rect 29920 21490 29972 21496
rect 29736 21004 29788 21010
rect 29736 20946 29788 20952
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29644 19372 29696 19378
rect 29644 19314 29696 19320
rect 28816 18964 28868 18970
rect 28816 18906 28868 18912
rect 28724 18692 28776 18698
rect 28724 18634 28776 18640
rect 28736 18578 28764 18634
rect 28736 18550 28856 18578
rect 28828 18426 28856 18550
rect 28356 18420 28408 18426
rect 28356 18362 28408 18368
rect 28816 18420 28868 18426
rect 28816 18362 28868 18368
rect 28264 17808 28316 17814
rect 28264 17750 28316 17756
rect 28276 17338 28304 17750
rect 28828 17678 28856 18362
rect 29748 18290 29776 20946
rect 29932 19854 29960 21490
rect 30024 21010 30052 21966
rect 30300 21622 30328 22578
rect 30288 21616 30340 21622
rect 30288 21558 30340 21564
rect 30012 21004 30064 21010
rect 30012 20946 30064 20952
rect 29920 19848 29972 19854
rect 29920 19790 29972 19796
rect 29828 19168 29880 19174
rect 29828 19110 29880 19116
rect 29920 19168 29972 19174
rect 29920 19110 29972 19116
rect 29840 18290 29868 19110
rect 29736 18284 29788 18290
rect 29736 18226 29788 18232
rect 29828 18284 29880 18290
rect 29828 18226 29880 18232
rect 29748 17898 29776 18226
rect 29748 17882 29868 17898
rect 29748 17876 29880 17882
rect 29748 17870 29828 17876
rect 28816 17672 28868 17678
rect 28816 17614 28868 17620
rect 29000 17536 29052 17542
rect 29000 17478 29052 17484
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28724 17264 28776 17270
rect 28724 17206 28776 17212
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28460 16794 28488 17138
rect 28448 16788 28500 16794
rect 28448 16730 28500 16736
rect 28736 16114 28764 17206
rect 28908 16584 28960 16590
rect 29012 16574 29040 17478
rect 29748 17202 29776 17870
rect 29828 17818 29880 17824
rect 29736 17196 29788 17202
rect 29736 17138 29788 17144
rect 28960 16546 29040 16574
rect 28908 16526 28960 16532
rect 29092 16448 29144 16454
rect 29092 16390 29144 16396
rect 29104 16182 29132 16390
rect 29092 16176 29144 16182
rect 29092 16118 29144 16124
rect 28724 16108 28776 16114
rect 28724 16050 28776 16056
rect 28816 16108 28868 16114
rect 28816 16050 28868 16056
rect 28540 15496 28592 15502
rect 28538 15464 28540 15473
rect 28592 15464 28594 15473
rect 28538 15399 28594 15408
rect 28736 14958 28764 16050
rect 28828 15706 28856 16050
rect 29368 15904 29420 15910
rect 29368 15846 29420 15852
rect 28816 15700 28868 15706
rect 28816 15642 28868 15648
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 29104 15502 29132 15642
rect 29092 15496 29144 15502
rect 28906 15464 28962 15473
rect 29144 15444 29224 15450
rect 29092 15438 29224 15444
rect 29104 15422 29224 15438
rect 28906 15399 28962 15408
rect 28920 15366 28948 15399
rect 28908 15360 28960 15366
rect 28908 15302 28960 15308
rect 28908 15020 28960 15026
rect 28908 14962 28960 14968
rect 28724 14952 28776 14958
rect 28724 14894 28776 14900
rect 28080 14884 28132 14890
rect 28080 14826 28132 14832
rect 27986 14512 28042 14521
rect 27986 14447 28042 14456
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27528 14340 27580 14346
rect 27528 14282 27580 14288
rect 27712 14340 27764 14346
rect 27712 14282 27764 14288
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 14074 27936 14282
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 28000 13462 28028 14350
rect 28092 14006 28120 14826
rect 28736 14482 28764 14894
rect 28920 14822 28948 14962
rect 28908 14816 28960 14822
rect 28908 14758 28960 14764
rect 28724 14476 28776 14482
rect 28724 14418 28776 14424
rect 28080 14000 28132 14006
rect 28080 13942 28132 13948
rect 27344 13456 27396 13462
rect 27344 13398 27396 13404
rect 27988 13456 28040 13462
rect 27988 13398 28040 13404
rect 27436 13388 27488 13394
rect 27436 13330 27488 13336
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27448 12850 27476 13330
rect 28092 12918 28120 13942
rect 28736 13938 28764 14418
rect 28908 14340 28960 14346
rect 28908 14282 28960 14288
rect 28632 13932 28684 13938
rect 28632 13874 28684 13880
rect 28724 13932 28776 13938
rect 28724 13874 28776 13880
rect 28356 13728 28408 13734
rect 28356 13670 28408 13676
rect 28264 13252 28316 13258
rect 28264 13194 28316 13200
rect 28276 12986 28304 13194
rect 28264 12980 28316 12986
rect 28264 12922 28316 12928
rect 28080 12912 28132 12918
rect 28080 12854 28132 12860
rect 28368 12850 28396 13670
rect 28644 13326 28672 13874
rect 28920 13326 28948 14282
rect 29000 14272 29052 14278
rect 29000 14214 29052 14220
rect 29012 13462 29040 14214
rect 29196 14006 29224 15422
rect 29380 15366 29408 15846
rect 29368 15360 29420 15366
rect 29368 15302 29420 15308
rect 29380 15026 29408 15302
rect 29368 15020 29420 15026
rect 29368 14962 29420 14968
rect 29184 14000 29236 14006
rect 29184 13942 29236 13948
rect 29092 13932 29144 13938
rect 29092 13874 29144 13880
rect 29104 13530 29132 13874
rect 29092 13524 29144 13530
rect 29092 13466 29144 13472
rect 29000 13456 29052 13462
rect 29000 13398 29052 13404
rect 29196 13326 29224 13942
rect 28632 13320 28684 13326
rect 28632 13262 28684 13268
rect 28908 13320 28960 13326
rect 28908 13262 28960 13268
rect 29184 13320 29236 13326
rect 29184 13262 29236 13268
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 27436 12844 27488 12850
rect 27436 12786 27488 12792
rect 28356 12844 28408 12850
rect 28356 12786 28408 12792
rect 27252 12776 27304 12782
rect 27252 12718 27304 12724
rect 26792 12300 26844 12306
rect 26792 12242 26844 12248
rect 27264 12238 27292 12718
rect 27344 12436 27396 12442
rect 27448 12434 27476 12786
rect 27396 12406 27476 12434
rect 27344 12378 27396 12384
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 26700 12164 26752 12170
rect 26700 12106 26752 12112
rect 24032 11892 24084 11898
rect 24032 11834 24084 11840
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 20536 11552 20588 11558
rect 20536 11494 20588 11500
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19352 6886 19472 6914
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 1860 2508 1912 2514
rect 1860 2450 1912 2456
rect 19444 2446 19472 6886
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 29656 2650 29684 13262
rect 29932 8974 29960 19110
rect 30196 17196 30248 17202
rect 30196 17138 30248 17144
rect 30208 16794 30236 17138
rect 30196 16788 30248 16794
rect 30196 16730 30248 16736
rect 30208 16658 30236 16730
rect 30196 16652 30248 16658
rect 30196 16594 30248 16600
rect 30392 15706 30420 22630
rect 30564 22500 30616 22506
rect 30564 22442 30616 22448
rect 30576 20942 30604 22442
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30564 20936 30616 20942
rect 30564 20878 30616 20884
rect 30944 20398 30972 21286
rect 31128 20602 31156 22646
rect 31116 20596 31168 20602
rect 31116 20538 31168 20544
rect 30564 20392 30616 20398
rect 30564 20334 30616 20340
rect 30932 20392 30984 20398
rect 30932 20334 30984 20340
rect 30576 19854 30604 20334
rect 30564 19848 30616 19854
rect 30564 19790 30616 19796
rect 30472 19508 30524 19514
rect 30472 19450 30524 19456
rect 30484 17270 30512 19450
rect 30576 17678 30604 19790
rect 30932 19712 30984 19718
rect 30932 19654 30984 19660
rect 30944 19378 30972 19654
rect 30932 19372 30984 19378
rect 30932 19314 30984 19320
rect 31220 18766 31248 23258
rect 31772 23118 31800 24006
rect 31956 23526 31984 24686
rect 32048 24206 32076 26182
rect 32312 24812 32364 24818
rect 32312 24754 32364 24760
rect 32128 24608 32180 24614
rect 32128 24550 32180 24556
rect 32140 24206 32168 24550
rect 32036 24200 32088 24206
rect 32036 24142 32088 24148
rect 32128 24200 32180 24206
rect 32128 24142 32180 24148
rect 32048 23730 32076 24142
rect 32036 23724 32088 23730
rect 32036 23666 32088 23672
rect 31944 23520 31996 23526
rect 31944 23462 31996 23468
rect 31956 23186 31984 23462
rect 31944 23180 31996 23186
rect 31944 23122 31996 23128
rect 31760 23112 31812 23118
rect 31760 23054 31812 23060
rect 31484 22432 31536 22438
rect 31484 22374 31536 22380
rect 31496 22030 31524 22374
rect 31772 22234 31800 23054
rect 32048 22642 32076 23666
rect 32324 23254 32352 24754
rect 32600 24614 32628 26386
rect 32588 24608 32640 24614
rect 32588 24550 32640 24556
rect 32588 23520 32640 23526
rect 32588 23462 32640 23468
rect 32312 23248 32364 23254
rect 32312 23190 32364 23196
rect 32600 22710 32628 23462
rect 32588 22704 32640 22710
rect 32588 22646 32640 22652
rect 32036 22636 32088 22642
rect 32036 22578 32088 22584
rect 31760 22228 31812 22234
rect 31760 22170 31812 22176
rect 31484 22024 31536 22030
rect 31484 21966 31536 21972
rect 31392 21888 31444 21894
rect 31392 21830 31444 21836
rect 31404 21622 31432 21830
rect 31772 21690 31800 22170
rect 32496 22024 32548 22030
rect 32496 21966 32548 21972
rect 32588 22024 32640 22030
rect 32588 21966 32640 21972
rect 31760 21684 31812 21690
rect 31760 21626 31812 21632
rect 31392 21616 31444 21622
rect 31392 21558 31444 21564
rect 32404 20936 32456 20942
rect 32404 20878 32456 20884
rect 31668 20800 31720 20806
rect 31668 20742 31720 20748
rect 31680 20398 31708 20742
rect 31668 20392 31720 20398
rect 31668 20334 31720 20340
rect 31392 20256 31444 20262
rect 31392 20198 31444 20204
rect 31404 19310 31432 20198
rect 31680 19922 31708 20334
rect 31668 19916 31720 19922
rect 31668 19858 31720 19864
rect 32416 19854 32444 20878
rect 32508 20806 32536 21966
rect 32600 21690 32628 21966
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32588 21548 32640 21554
rect 32588 21490 32640 21496
rect 32496 20800 32548 20806
rect 32496 20742 32548 20748
rect 32508 20534 32536 20742
rect 32600 20602 32628 21490
rect 32680 21412 32732 21418
rect 32680 21354 32732 21360
rect 32588 20596 32640 20602
rect 32588 20538 32640 20544
rect 32496 20528 32548 20534
rect 32496 20470 32548 20476
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 32404 19848 32456 19854
rect 32404 19790 32456 19796
rect 31588 19378 31616 19790
rect 31576 19372 31628 19378
rect 31576 19314 31628 19320
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 31392 19304 31444 19310
rect 31392 19246 31444 19252
rect 31208 18760 31260 18766
rect 31208 18702 31260 18708
rect 31220 18154 31248 18702
rect 31208 18148 31260 18154
rect 31208 18090 31260 18096
rect 31220 17678 31248 18090
rect 30564 17672 30616 17678
rect 30564 17614 30616 17620
rect 31208 17672 31260 17678
rect 31208 17614 31260 17620
rect 30748 17536 30800 17542
rect 30748 17478 30800 17484
rect 30472 17264 30524 17270
rect 30472 17206 30524 17212
rect 30564 16516 30616 16522
rect 30564 16458 30616 16464
rect 30576 16250 30604 16458
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30760 16114 30788 17478
rect 30840 16516 30892 16522
rect 30840 16458 30892 16464
rect 30748 16108 30800 16114
rect 30748 16050 30800 16056
rect 30852 15706 30880 16458
rect 30932 15904 30984 15910
rect 30932 15846 30984 15852
rect 30380 15700 30432 15706
rect 30380 15642 30432 15648
rect 30840 15700 30892 15706
rect 30840 15642 30892 15648
rect 30944 15502 30972 15846
rect 30932 15496 30984 15502
rect 30932 15438 30984 15444
rect 30656 15360 30708 15366
rect 30656 15302 30708 15308
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30024 14618 30052 14962
rect 30012 14612 30064 14618
rect 30012 14554 30064 14560
rect 30668 14414 30696 15302
rect 31404 15162 31432 19246
rect 32324 17678 32352 19314
rect 32416 18834 32444 19790
rect 32692 19514 32720 21354
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32588 19372 32640 19378
rect 32588 19314 32640 19320
rect 32496 19168 32548 19174
rect 32496 19110 32548 19116
rect 32404 18828 32456 18834
rect 32404 18770 32456 18776
rect 32416 18290 32444 18770
rect 32404 18284 32456 18290
rect 32404 18226 32456 18232
rect 32508 17746 32536 19110
rect 32496 17740 32548 17746
rect 32496 17682 32548 17688
rect 32312 17672 32364 17678
rect 32312 17614 32364 17620
rect 31576 17604 31628 17610
rect 31576 17546 31628 17552
rect 31588 16114 31616 17546
rect 32220 17264 32272 17270
rect 32220 17206 32272 17212
rect 32232 16574 32260 17206
rect 32324 17134 32352 17614
rect 32508 17270 32536 17682
rect 32600 17338 32628 19314
rect 32588 17332 32640 17338
rect 32588 17274 32640 17280
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32508 17066 32536 17206
rect 32496 17060 32548 17066
rect 32496 17002 32548 17008
rect 32140 16546 32260 16574
rect 32140 16454 32168 16546
rect 32128 16448 32180 16454
rect 32128 16390 32180 16396
rect 31576 16108 31628 16114
rect 31576 16050 31628 16056
rect 32140 16046 32168 16390
rect 32128 16040 32180 16046
rect 32128 15982 32180 15988
rect 31484 15972 31536 15978
rect 31484 15914 31536 15920
rect 31496 15502 31524 15914
rect 32680 15904 32732 15910
rect 32680 15846 32732 15852
rect 31484 15496 31536 15502
rect 31484 15438 31536 15444
rect 31392 15156 31444 15162
rect 31392 15098 31444 15104
rect 32588 14952 32640 14958
rect 32588 14894 32640 14900
rect 32600 14618 32628 14894
rect 32692 14822 32720 15846
rect 32680 14816 32732 14822
rect 32680 14758 32732 14764
rect 32588 14612 32640 14618
rect 32588 14554 32640 14560
rect 30196 14408 30248 14414
rect 30196 14350 30248 14356
rect 30656 14408 30708 14414
rect 30656 14350 30708 14356
rect 30208 13530 30236 14350
rect 30196 13524 30248 13530
rect 30196 13466 30248 13472
rect 32784 13394 32812 27066
rect 32876 27062 32904 29106
rect 33520 29034 33548 29124
rect 33416 29028 33468 29034
rect 33416 28970 33468 28976
rect 33508 29028 33560 29034
rect 33508 28970 33560 28976
rect 33428 28558 33456 28970
rect 33416 28552 33468 28558
rect 33416 28494 33468 28500
rect 33232 28416 33284 28422
rect 33232 28358 33284 28364
rect 33244 28150 33272 28358
rect 33232 28144 33284 28150
rect 33232 28086 33284 28092
rect 33704 27606 33732 30262
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 33980 28966 34008 29582
rect 33968 28960 34020 28966
rect 33968 28902 34020 28908
rect 33324 27600 33376 27606
rect 33324 27542 33376 27548
rect 33692 27600 33744 27606
rect 33692 27542 33744 27548
rect 32864 27056 32916 27062
rect 32864 26998 32916 27004
rect 33336 26518 33364 27542
rect 33600 27532 33652 27538
rect 33600 27474 33652 27480
rect 33612 26994 33640 27474
rect 34072 27470 34100 30534
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34164 29850 34192 30194
rect 34152 29844 34204 29850
rect 34152 29786 34204 29792
rect 34244 29572 34296 29578
rect 34244 29514 34296 29520
rect 34152 29504 34204 29510
rect 34152 29446 34204 29452
rect 34164 29238 34192 29446
rect 34256 29306 34284 29514
rect 34244 29300 34296 29306
rect 34244 29242 34296 29248
rect 34152 29232 34204 29238
rect 34152 29174 34204 29180
rect 34336 29232 34388 29238
rect 34336 29174 34388 29180
rect 34164 28626 34192 29174
rect 34152 28620 34204 28626
rect 34152 28562 34204 28568
rect 34164 28218 34192 28562
rect 34348 28558 34376 29174
rect 34336 28552 34388 28558
rect 34336 28494 34388 28500
rect 34152 28212 34204 28218
rect 34152 28154 34204 28160
rect 34336 28076 34388 28082
rect 34336 28018 34388 28024
rect 34348 27674 34376 28018
rect 34336 27668 34388 27674
rect 34336 27610 34388 27616
rect 34060 27464 34112 27470
rect 34060 27406 34112 27412
rect 34060 27328 34112 27334
rect 34060 27270 34112 27276
rect 33600 26988 33652 26994
rect 33600 26930 33652 26936
rect 33324 26512 33376 26518
rect 33324 26454 33376 26460
rect 33336 25498 33364 26454
rect 33612 26382 33640 26930
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 33612 26234 33640 26318
rect 33692 26308 33744 26314
rect 33692 26250 33744 26256
rect 33428 26206 33640 26234
rect 33324 25492 33376 25498
rect 33324 25434 33376 25440
rect 33428 25378 33456 26206
rect 33508 25492 33560 25498
rect 33508 25434 33560 25440
rect 33336 25350 33456 25378
rect 33336 25226 33364 25350
rect 32956 25220 33008 25226
rect 32956 25162 33008 25168
rect 33324 25220 33376 25226
rect 33324 25162 33376 25168
rect 32968 24682 32996 25162
rect 32956 24676 33008 24682
rect 32956 24618 33008 24624
rect 32864 23860 32916 23866
rect 32864 23802 32916 23808
rect 32876 23254 32904 23802
rect 32968 23798 32996 24618
rect 33048 24608 33100 24614
rect 33048 24550 33100 24556
rect 32956 23792 33008 23798
rect 32956 23734 33008 23740
rect 32864 23248 32916 23254
rect 32864 23190 32916 23196
rect 33060 23118 33088 24550
rect 33048 23112 33100 23118
rect 33048 23054 33100 23060
rect 33140 23078 33192 23084
rect 33140 23020 33192 23026
rect 33152 22642 33180 23020
rect 33140 22636 33192 22642
rect 33140 22578 33192 22584
rect 33336 22420 33364 25162
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 33428 24410 33456 24686
rect 33416 24404 33468 24410
rect 33416 24346 33468 24352
rect 33428 23662 33456 24346
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 33520 23118 33548 25434
rect 33704 24818 33732 26250
rect 34072 25498 34100 27270
rect 34440 26042 34468 31214
rect 34624 30190 34652 31758
rect 35544 31346 35572 31758
rect 36728 31680 36780 31686
rect 36728 31622 36780 31628
rect 36740 31414 36768 31622
rect 36728 31408 36780 31414
rect 36728 31350 36780 31356
rect 35532 31340 35584 31346
rect 35532 31282 35584 31288
rect 36176 31340 36228 31346
rect 36176 31282 36228 31288
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35544 30870 35572 31282
rect 36188 30938 36216 31282
rect 36924 30938 36952 31758
rect 36176 30932 36228 30938
rect 36176 30874 36228 30880
rect 36912 30932 36964 30938
rect 36912 30874 36964 30880
rect 35532 30864 35584 30870
rect 35532 30806 35584 30812
rect 35544 30394 35572 30806
rect 36188 30734 36216 30874
rect 36912 30796 36964 30802
rect 36912 30738 36964 30744
rect 35716 30728 35768 30734
rect 35716 30670 35768 30676
rect 36176 30728 36228 30734
rect 36176 30670 36228 30676
rect 35624 30592 35676 30598
rect 35624 30534 35676 30540
rect 35532 30388 35584 30394
rect 35532 30330 35584 30336
rect 35636 30326 35664 30534
rect 35624 30320 35676 30326
rect 35624 30262 35676 30268
rect 34796 30252 34848 30258
rect 34796 30194 34848 30200
rect 34612 30184 34664 30190
rect 34612 30126 34664 30132
rect 34520 29640 34572 29646
rect 34520 29582 34572 29588
rect 34532 29102 34560 29582
rect 34520 29096 34572 29102
rect 34520 29038 34572 29044
rect 34624 27946 34652 30126
rect 34808 29850 34836 30194
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29844 34848 29850
rect 34796 29786 34848 29792
rect 35728 29306 35756 30670
rect 36268 30660 36320 30666
rect 36268 30602 36320 30608
rect 36280 30326 36308 30602
rect 36268 30320 36320 30326
rect 36268 30262 36320 30268
rect 36280 29850 36308 30262
rect 36268 29844 36320 29850
rect 36268 29786 36320 29792
rect 36924 29714 36952 30738
rect 37200 30734 37228 32166
rect 37280 31952 37332 31958
rect 37280 31894 37332 31900
rect 37188 30728 37240 30734
rect 37188 30670 37240 30676
rect 36912 29708 36964 29714
rect 36912 29650 36964 29656
rect 35992 29572 36044 29578
rect 35992 29514 36044 29520
rect 35716 29300 35768 29306
rect 35716 29242 35768 29248
rect 36004 29238 36032 29514
rect 35992 29232 36044 29238
rect 35992 29174 36044 29180
rect 35348 29164 35400 29170
rect 35348 29106 35400 29112
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34796 28484 34848 28490
rect 34796 28426 34848 28432
rect 34808 28218 34836 28426
rect 35360 28422 35388 29106
rect 36176 28960 36228 28966
rect 36176 28902 36228 28908
rect 35532 28756 35584 28762
rect 35532 28698 35584 28704
rect 34980 28416 35032 28422
rect 34980 28358 35032 28364
rect 35348 28416 35400 28422
rect 35348 28358 35400 28364
rect 34796 28212 34848 28218
rect 34796 28154 34848 28160
rect 34992 28082 35020 28358
rect 34980 28076 35032 28082
rect 34980 28018 35032 28024
rect 34612 27940 34664 27946
rect 34612 27882 34664 27888
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35544 27674 35572 28698
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 36004 28218 36032 28426
rect 35992 28212 36044 28218
rect 35992 28154 36044 28160
rect 36188 28082 36216 28902
rect 36924 28642 36952 29650
rect 37292 29170 37320 31894
rect 37464 31680 37516 31686
rect 37464 31622 37516 31628
rect 37372 31136 37424 31142
rect 37372 31078 37424 31084
rect 37384 30122 37412 31078
rect 37372 30116 37424 30122
rect 37372 30058 37424 30064
rect 37384 29578 37412 30058
rect 37476 29646 37504 31622
rect 37660 31482 37688 32370
rect 37832 31816 37884 31822
rect 37832 31758 37884 31764
rect 38292 31816 38344 31822
rect 38292 31758 38344 31764
rect 37648 31476 37700 31482
rect 37648 31418 37700 31424
rect 37556 30252 37608 30258
rect 37556 30194 37608 30200
rect 37568 29850 37596 30194
rect 37556 29844 37608 29850
rect 37556 29786 37608 29792
rect 37464 29640 37516 29646
rect 37464 29582 37516 29588
rect 37372 29572 37424 29578
rect 37372 29514 37424 29520
rect 37844 29306 37872 31758
rect 37924 30592 37976 30598
rect 37924 30534 37976 30540
rect 37936 30394 37964 30534
rect 37924 30388 37976 30394
rect 37924 30330 37976 30336
rect 37832 29300 37884 29306
rect 37832 29242 37884 29248
rect 37936 29238 37964 30330
rect 38304 29345 38332 31758
rect 38290 29336 38346 29345
rect 38290 29271 38346 29280
rect 37924 29232 37976 29238
rect 37924 29174 37976 29180
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37648 29164 37700 29170
rect 37648 29106 37700 29112
rect 36832 28614 36952 28642
rect 36832 28558 36860 28614
rect 36820 28552 36872 28558
rect 36820 28494 36872 28500
rect 36176 28076 36228 28082
rect 36176 28018 36228 28024
rect 36728 27872 36780 27878
rect 36728 27814 36780 27820
rect 35532 27668 35584 27674
rect 35532 27610 35584 27616
rect 35072 27464 35124 27470
rect 35072 27406 35124 27412
rect 35084 27130 35112 27406
rect 35348 27328 35400 27334
rect 35348 27270 35400 27276
rect 35072 27124 35124 27130
rect 35072 27066 35124 27072
rect 35360 26994 35388 27270
rect 35348 26988 35400 26994
rect 35348 26930 35400 26936
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34612 26512 34664 26518
rect 34612 26454 34664 26460
rect 34624 26314 34652 26454
rect 35360 26450 35388 26930
rect 35544 26790 35572 27610
rect 36740 27470 36768 27814
rect 36832 27674 36860 28494
rect 37660 28082 37688 29106
rect 37556 28076 37608 28082
rect 37556 28018 37608 28024
rect 37648 28076 37700 28082
rect 37648 28018 37700 28024
rect 37464 27872 37516 27878
rect 37464 27814 37516 27820
rect 36820 27668 36872 27674
rect 36820 27610 36872 27616
rect 35624 27464 35676 27470
rect 35624 27406 35676 27412
rect 35808 27464 35860 27470
rect 35808 27406 35860 27412
rect 36728 27464 36780 27470
rect 36728 27406 36780 27412
rect 35532 26784 35584 26790
rect 35532 26726 35584 26732
rect 35348 26444 35400 26450
rect 35348 26386 35400 26392
rect 35636 26382 35664 27406
rect 35820 27130 35848 27406
rect 36452 27328 36504 27334
rect 36452 27270 36504 27276
rect 35808 27124 35860 27130
rect 35808 27066 35860 27072
rect 35256 26376 35308 26382
rect 35256 26318 35308 26324
rect 35624 26376 35676 26382
rect 35624 26318 35676 26324
rect 34612 26308 34664 26314
rect 34612 26250 34664 26256
rect 34428 26036 34480 26042
rect 34428 25978 34480 25984
rect 34520 25968 34572 25974
rect 34520 25910 34572 25916
rect 34060 25492 34112 25498
rect 34060 25434 34112 25440
rect 34532 25294 34560 25910
rect 34520 25288 34572 25294
rect 34520 25230 34572 25236
rect 33876 25152 33928 25158
rect 33876 25094 33928 25100
rect 33888 24886 33916 25094
rect 33876 24880 33928 24886
rect 33876 24822 33928 24828
rect 33692 24812 33744 24818
rect 33692 24754 33744 24760
rect 33888 24138 33916 24822
rect 33876 24132 33928 24138
rect 33876 24074 33928 24080
rect 33784 23724 33836 23730
rect 33784 23666 33836 23672
rect 33796 23322 33824 23666
rect 33784 23316 33836 23322
rect 33784 23258 33836 23264
rect 33508 23112 33560 23118
rect 33508 23054 33560 23060
rect 33416 22432 33468 22438
rect 33336 22392 33416 22420
rect 33416 22374 33468 22380
rect 33140 22092 33192 22098
rect 33140 22034 33192 22040
rect 33152 20874 33180 22034
rect 33140 20868 33192 20874
rect 33140 20810 33192 20816
rect 33152 20602 33180 20810
rect 33140 20596 33192 20602
rect 33140 20538 33192 20544
rect 33428 20448 33456 22374
rect 33520 21962 33548 23054
rect 33888 23050 33916 24074
rect 34244 23588 34296 23594
rect 34244 23530 34296 23536
rect 34256 23322 34284 23530
rect 34244 23316 34296 23322
rect 34244 23258 34296 23264
rect 33692 23044 33744 23050
rect 33692 22986 33744 22992
rect 33876 23044 33928 23050
rect 33876 22986 33928 22992
rect 34520 23044 34572 23050
rect 34520 22986 34572 22992
rect 33704 22778 33732 22986
rect 33692 22772 33744 22778
rect 33692 22714 33744 22720
rect 33968 22772 34020 22778
rect 33968 22714 34020 22720
rect 33600 22024 33652 22030
rect 33600 21966 33652 21972
rect 33508 21956 33560 21962
rect 33508 21898 33560 21904
rect 33520 21622 33548 21898
rect 33508 21616 33560 21622
rect 33508 21558 33560 21564
rect 33508 20460 33560 20466
rect 33428 20420 33508 20448
rect 33508 20402 33560 20408
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 20256 33192 20262
rect 33140 20198 33192 20204
rect 33152 19530 33180 20198
rect 33244 20058 33272 20334
rect 33324 20324 33376 20330
rect 33324 20266 33376 20272
rect 33232 20052 33284 20058
rect 33232 19994 33284 20000
rect 32864 19508 32916 19514
rect 33152 19502 33272 19530
rect 32864 19450 32916 19456
rect 32876 17338 32904 19450
rect 33244 19446 33272 19502
rect 33140 19440 33192 19446
rect 33140 19382 33192 19388
rect 33232 19440 33284 19446
rect 33232 19382 33284 19388
rect 33152 18766 33180 19382
rect 33232 19304 33284 19310
rect 33232 19246 33284 19252
rect 33140 18760 33192 18766
rect 33140 18702 33192 18708
rect 33244 18426 33272 19246
rect 33336 19174 33364 20266
rect 33520 19922 33548 20402
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33416 19780 33468 19786
rect 33416 19722 33468 19728
rect 33324 19168 33376 19174
rect 33324 19110 33376 19116
rect 33428 18970 33456 19722
rect 33612 19514 33640 21966
rect 33600 19508 33652 19514
rect 33600 19450 33652 19456
rect 33416 18964 33468 18970
rect 33416 18906 33468 18912
rect 33232 18420 33284 18426
rect 33232 18362 33284 18368
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 33244 17270 33272 18362
rect 33416 17672 33468 17678
rect 33416 17614 33468 17620
rect 33232 17264 33284 17270
rect 33232 17206 33284 17212
rect 33428 16794 33456 17614
rect 33416 16788 33468 16794
rect 33416 16730 33468 16736
rect 33980 16726 34008 22714
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 34440 22234 34468 22578
rect 34428 22228 34480 22234
rect 34428 22170 34480 22176
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 34164 21486 34192 21966
rect 34152 21480 34204 21486
rect 34152 21422 34204 21428
rect 34532 19281 34560 22986
rect 34518 19272 34574 19281
rect 34518 19207 34574 19216
rect 34244 18760 34296 18766
rect 34244 18702 34296 18708
rect 34520 18760 34572 18766
rect 34520 18702 34572 18708
rect 34060 18624 34112 18630
rect 34060 18566 34112 18572
rect 34072 18358 34100 18566
rect 34060 18352 34112 18358
rect 34060 18294 34112 18300
rect 34256 17882 34284 18702
rect 34428 18080 34480 18086
rect 34428 18022 34480 18028
rect 34244 17876 34296 17882
rect 34244 17818 34296 17824
rect 34440 17270 34468 18022
rect 34428 17264 34480 17270
rect 34428 17206 34480 17212
rect 34532 16998 34560 18702
rect 34624 18170 34652 26250
rect 34888 26240 34940 26246
rect 34888 26182 34940 26188
rect 34796 25968 34848 25974
rect 34796 25910 34848 25916
rect 34808 25838 34836 25910
rect 34900 25906 34928 26182
rect 35268 25974 35296 26318
rect 35820 26314 35848 27066
rect 36464 26994 36492 27270
rect 36832 27062 36860 27610
rect 36820 27056 36872 27062
rect 36820 26998 36872 27004
rect 36360 26988 36412 26994
rect 36360 26930 36412 26936
rect 36452 26988 36504 26994
rect 36452 26930 36504 26936
rect 36636 26988 36688 26994
rect 36636 26930 36688 26936
rect 36176 26784 36228 26790
rect 36176 26726 36228 26732
rect 36188 26450 36216 26726
rect 36372 26586 36400 26930
rect 36360 26580 36412 26586
rect 36360 26522 36412 26528
rect 36176 26444 36228 26450
rect 36176 26386 36228 26392
rect 35808 26308 35860 26314
rect 35808 26250 35860 26256
rect 36176 26308 36228 26314
rect 36176 26250 36228 26256
rect 36188 26042 36216 26250
rect 36176 26036 36228 26042
rect 36176 25978 36228 25984
rect 35256 25968 35308 25974
rect 35256 25910 35308 25916
rect 34888 25900 34940 25906
rect 34888 25842 34940 25848
rect 36648 25838 36676 26930
rect 36832 26450 36860 26998
rect 36912 26852 36964 26858
rect 36912 26794 36964 26800
rect 36820 26444 36872 26450
rect 36820 26386 36872 26392
rect 36832 26234 36860 26386
rect 36740 26206 36860 26234
rect 34796 25832 34848 25838
rect 34796 25774 34848 25780
rect 36636 25832 36688 25838
rect 36636 25774 36688 25780
rect 35348 25696 35400 25702
rect 35348 25638 35400 25644
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34980 25220 35032 25226
rect 34980 25162 35032 25168
rect 34992 24954 35020 25162
rect 34980 24948 35032 24954
rect 34980 24890 35032 24896
rect 35360 24818 35388 25638
rect 36740 25362 36768 26206
rect 36728 25356 36780 25362
rect 36728 25298 36780 25304
rect 36176 25288 36228 25294
rect 36176 25230 36228 25236
rect 35348 24812 35400 24818
rect 35348 24754 35400 24760
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 36188 24274 36216 25230
rect 36924 24682 36952 26794
rect 37280 26240 37332 26246
rect 37280 26182 37332 26188
rect 37188 25832 37240 25838
rect 37188 25774 37240 25780
rect 37004 25696 37056 25702
rect 37004 25638 37056 25644
rect 37016 25294 37044 25638
rect 37004 25288 37056 25294
rect 37004 25230 37056 25236
rect 37200 25158 37228 25774
rect 37188 25152 37240 25158
rect 37188 25094 37240 25100
rect 37200 24954 37228 25094
rect 37188 24948 37240 24954
rect 37188 24890 37240 24896
rect 36912 24676 36964 24682
rect 36912 24618 36964 24624
rect 37200 24614 37228 24890
rect 37292 24682 37320 26182
rect 37476 26042 37504 27814
rect 37568 27130 37596 28018
rect 37556 27124 37608 27130
rect 37556 27066 37608 27072
rect 37660 26994 37688 28018
rect 38016 28008 38068 28014
rect 38016 27950 38068 27956
rect 38028 27334 38056 27950
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 37464 26036 37516 26042
rect 37464 25978 37516 25984
rect 37660 25906 37688 26930
rect 38028 26926 38056 27270
rect 38016 26920 38068 26926
rect 38016 26862 38068 26868
rect 37648 25900 37700 25906
rect 37648 25842 37700 25848
rect 37648 25152 37700 25158
rect 37648 25094 37700 25100
rect 37660 24818 37688 25094
rect 38292 24880 38344 24886
rect 38292 24822 38344 24828
rect 37464 24812 37516 24818
rect 37464 24754 37516 24760
rect 37648 24812 37700 24818
rect 37648 24754 37700 24760
rect 37280 24676 37332 24682
rect 37280 24618 37332 24624
rect 37188 24608 37240 24614
rect 37188 24550 37240 24556
rect 36176 24268 36228 24274
rect 36176 24210 36228 24216
rect 34796 24064 34848 24070
rect 34796 24006 34848 24012
rect 34808 23050 34836 24006
rect 36188 23798 36216 24210
rect 36636 24132 36688 24138
rect 36636 24074 36688 24080
rect 36648 23866 36676 24074
rect 36636 23860 36688 23866
rect 36636 23802 36688 23808
rect 35532 23792 35584 23798
rect 35532 23734 35584 23740
rect 36176 23792 36228 23798
rect 36176 23734 36228 23740
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35544 23118 35572 23734
rect 36188 23186 36216 23734
rect 37476 23730 37504 24754
rect 37556 24744 37608 24750
rect 37556 24686 37608 24692
rect 37568 24410 37596 24686
rect 37556 24404 37608 24410
rect 37556 24346 37608 24352
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37648 23724 37700 23730
rect 37648 23666 37700 23672
rect 36176 23180 36228 23186
rect 36176 23122 36228 23128
rect 34888 23112 34940 23118
rect 34888 23054 34940 23060
rect 35532 23112 35584 23118
rect 35532 23054 35584 23060
rect 34796 23044 34848 23050
rect 34796 22986 34848 22992
rect 34900 22642 34928 23054
rect 35532 22976 35584 22982
rect 35532 22918 35584 22924
rect 35808 22976 35860 22982
rect 35808 22918 35860 22924
rect 34888 22636 34940 22642
rect 34888 22578 34940 22584
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35164 22228 35216 22234
rect 35164 22170 35216 22176
rect 34704 22092 34756 22098
rect 34704 22034 34756 22040
rect 34716 21622 34744 22034
rect 35176 21962 35204 22170
rect 35544 22098 35572 22918
rect 35624 22432 35676 22438
rect 35624 22374 35676 22380
rect 35532 22092 35584 22098
rect 35532 22034 35584 22040
rect 35164 21956 35216 21962
rect 35164 21898 35216 21904
rect 35636 21894 35664 22374
rect 35820 22234 35848 22918
rect 37292 22778 37320 23666
rect 37556 23520 37608 23526
rect 37556 23462 37608 23468
rect 37372 23044 37424 23050
rect 37372 22986 37424 22992
rect 37280 22772 37332 22778
rect 37280 22714 37332 22720
rect 36268 22432 36320 22438
rect 36268 22374 36320 22380
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 36176 22092 36228 22098
rect 36176 22034 36228 22040
rect 35900 22024 35952 22030
rect 36188 21978 36216 22034
rect 36280 22030 36308 22374
rect 37384 22234 37412 22986
rect 37372 22228 37424 22234
rect 37372 22170 37424 22176
rect 37568 22030 37596 23462
rect 37660 22642 37688 23666
rect 38304 23322 38332 24822
rect 38292 23316 38344 23322
rect 38292 23258 38344 23264
rect 38304 22710 38332 23258
rect 38292 22704 38344 22710
rect 38292 22646 38344 22652
rect 37648 22636 37700 22642
rect 37648 22578 37700 22584
rect 35952 21972 36216 21978
rect 35900 21966 36216 21972
rect 36268 22024 36320 22030
rect 36268 21966 36320 21972
rect 37556 22024 37608 22030
rect 37556 21966 37608 21972
rect 35912 21950 36216 21966
rect 35348 21888 35400 21894
rect 35348 21830 35400 21836
rect 35624 21888 35676 21894
rect 35624 21830 35676 21836
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 34796 21480 34848 21486
rect 34796 21422 34848 21428
rect 34808 20534 34836 21422
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35360 21162 35388 21830
rect 36188 21690 36216 21950
rect 35716 21684 35768 21690
rect 35716 21626 35768 21632
rect 36176 21684 36228 21690
rect 36176 21626 36228 21632
rect 35624 21616 35676 21622
rect 35624 21558 35676 21564
rect 35636 21350 35664 21558
rect 35532 21344 35584 21350
rect 35532 21286 35584 21292
rect 35624 21344 35676 21350
rect 35624 21286 35676 21292
rect 35268 21134 35388 21162
rect 35268 20806 35296 21134
rect 35544 20942 35572 21286
rect 35532 20936 35584 20942
rect 35532 20878 35584 20884
rect 35256 20800 35308 20806
rect 35256 20742 35308 20748
rect 34796 20528 34848 20534
rect 34796 20470 34848 20476
rect 35268 20466 35296 20742
rect 35256 20460 35308 20466
rect 35256 20402 35308 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34704 19712 34756 19718
rect 34704 19654 34756 19660
rect 34716 19378 34744 19654
rect 34704 19372 34756 19378
rect 34704 19314 34756 19320
rect 35544 19310 35572 20878
rect 35728 19334 35756 21626
rect 37660 21622 37688 22578
rect 37648 21616 37700 21622
rect 37648 21558 37700 21564
rect 36636 21548 36688 21554
rect 36636 21490 36688 21496
rect 36176 21344 36228 21350
rect 36176 21286 36228 21292
rect 35992 20868 36044 20874
rect 35992 20810 36044 20816
rect 36004 20602 36032 20810
rect 35992 20596 36044 20602
rect 35992 20538 36044 20544
rect 36188 20466 36216 21286
rect 36648 20602 36676 21490
rect 36636 20596 36688 20602
rect 36636 20538 36688 20544
rect 36176 20460 36228 20466
rect 36176 20402 36228 20408
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 35808 19712 35860 19718
rect 35808 19654 35860 19660
rect 35820 19446 35848 19654
rect 35808 19440 35860 19446
rect 35808 19382 35860 19388
rect 35532 19304 35584 19310
rect 35728 19306 35940 19334
rect 35532 19246 35584 19252
rect 34704 19168 34756 19174
rect 34704 19110 34756 19116
rect 34716 18698 34744 19110
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35544 18766 35572 19246
rect 35532 18760 35584 18766
rect 35532 18702 35584 18708
rect 34704 18692 34756 18698
rect 34704 18634 34756 18640
rect 34716 18358 34744 18634
rect 34704 18352 34756 18358
rect 34704 18294 34756 18300
rect 35912 18290 35940 19306
rect 36004 18426 36032 19790
rect 36544 19780 36596 19786
rect 36544 19722 36596 19728
rect 36268 18624 36320 18630
rect 36268 18566 36320 18572
rect 35992 18420 36044 18426
rect 35992 18362 36044 18368
rect 36280 18358 36308 18566
rect 36268 18352 36320 18358
rect 36268 18294 36320 18300
rect 35900 18284 35952 18290
rect 35900 18226 35952 18232
rect 34704 18216 34756 18222
rect 34624 18164 34704 18170
rect 34624 18158 34756 18164
rect 35348 18216 35400 18222
rect 35348 18158 35400 18164
rect 34624 18142 34744 18158
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35360 17882 35388 18158
rect 35348 17876 35400 17882
rect 35348 17818 35400 17824
rect 35532 17672 35584 17678
rect 35532 17614 35584 17620
rect 34796 17604 34848 17610
rect 34796 17546 34848 17552
rect 34808 17338 34836 17546
rect 35544 17338 35572 17614
rect 35912 17610 35940 18226
rect 36556 18086 36584 19722
rect 37004 19508 37056 19514
rect 37004 19450 37056 19456
rect 36636 19168 36688 19174
rect 36636 19110 36688 19116
rect 36648 18170 36676 19110
rect 37016 18766 37044 19450
rect 37648 19372 37700 19378
rect 37648 19314 37700 19320
rect 37004 18760 37056 18766
rect 37004 18702 37056 18708
rect 37464 18624 37516 18630
rect 37464 18566 37516 18572
rect 37476 18222 37504 18566
rect 37556 18352 37608 18358
rect 37556 18294 37608 18300
rect 37464 18216 37516 18222
rect 36648 18142 36952 18170
rect 37464 18158 37516 18164
rect 36544 18080 36596 18086
rect 36544 18022 36596 18028
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 34796 17332 34848 17338
rect 34796 17274 34848 17280
rect 35532 17332 35584 17338
rect 35532 17274 35584 17280
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34532 16794 34560 16934
rect 34520 16788 34572 16794
rect 34520 16730 34572 16736
rect 33968 16720 34020 16726
rect 33968 16662 34020 16668
rect 33232 16244 33284 16250
rect 33232 16186 33284 16192
rect 32864 16108 32916 16114
rect 32916 16068 32996 16096
rect 32864 16050 32916 16056
rect 32968 15484 32996 16068
rect 33140 15904 33192 15910
rect 33140 15846 33192 15852
rect 33152 15570 33180 15846
rect 33244 15706 33272 16186
rect 33324 16108 33376 16114
rect 33324 16050 33376 16056
rect 33232 15700 33284 15706
rect 33232 15642 33284 15648
rect 33336 15570 33364 16050
rect 33980 16046 34008 16662
rect 34808 16590 34836 17274
rect 35440 17196 35492 17202
rect 35440 17138 35492 17144
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 34796 16584 34848 16590
rect 34796 16526 34848 16532
rect 34336 16448 34388 16454
rect 34336 16390 34388 16396
rect 34348 16114 34376 16390
rect 34336 16108 34388 16114
rect 34336 16050 34388 16056
rect 33968 16040 34020 16046
rect 33968 15982 34020 15988
rect 34808 15978 34836 16526
rect 35360 16522 35388 16934
rect 35348 16516 35400 16522
rect 35348 16458 35400 16464
rect 35452 16250 35480 17138
rect 35440 16244 35492 16250
rect 35440 16186 35492 16192
rect 35912 16114 35940 17546
rect 36556 17490 36584 18022
rect 36648 17678 36676 18142
rect 36924 18086 36952 18142
rect 36820 18080 36872 18086
rect 36820 18022 36872 18028
rect 36912 18080 36964 18086
rect 36912 18022 36964 18028
rect 36832 17814 36860 18022
rect 36820 17808 36872 17814
rect 36820 17750 36872 17756
rect 37476 17678 37504 18158
rect 36636 17672 36688 17678
rect 36636 17614 36688 17620
rect 37464 17672 37516 17678
rect 37464 17614 37516 17620
rect 36556 17462 36676 17490
rect 36268 17128 36320 17134
rect 36268 17070 36320 17076
rect 36280 16726 36308 17070
rect 36360 17060 36412 17066
rect 36360 17002 36412 17008
rect 36268 16720 36320 16726
rect 36268 16662 36320 16668
rect 36280 16250 36308 16662
rect 36268 16244 36320 16250
rect 36268 16186 36320 16192
rect 35900 16108 35952 16114
rect 35900 16050 35952 16056
rect 34796 15972 34848 15978
rect 34796 15914 34848 15920
rect 34808 15570 34836 15914
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35912 15638 35940 16050
rect 36372 15978 36400 17002
rect 36544 16992 36596 16998
rect 36544 16934 36596 16940
rect 36556 16182 36584 16934
rect 36544 16176 36596 16182
rect 36544 16118 36596 16124
rect 36176 15972 36228 15978
rect 36176 15914 36228 15920
rect 36360 15972 36412 15978
rect 36360 15914 36412 15920
rect 36188 15706 36216 15914
rect 36176 15700 36228 15706
rect 36176 15642 36228 15648
rect 35900 15632 35952 15638
rect 35900 15574 35952 15580
rect 33140 15564 33192 15570
rect 33140 15506 33192 15512
rect 33324 15564 33376 15570
rect 33324 15506 33376 15512
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 33048 15496 33100 15502
rect 32968 15456 33048 15484
rect 32968 14618 32996 15456
rect 33048 15438 33100 15444
rect 33152 15162 33180 15506
rect 36188 15502 36216 15642
rect 36176 15496 36228 15502
rect 36176 15438 36228 15444
rect 34888 15360 34940 15366
rect 34888 15302 34940 15308
rect 33140 15156 33192 15162
rect 33140 15098 33192 15104
rect 34900 15026 34928 15302
rect 36648 15162 36676 17462
rect 37280 17264 37332 17270
rect 37280 17206 37332 17212
rect 37188 16992 37240 16998
rect 37188 16934 37240 16940
rect 36912 16652 36964 16658
rect 36912 16594 36964 16600
rect 36924 15570 36952 16594
rect 37200 16590 37228 16934
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 37188 16448 37240 16454
rect 37188 16390 37240 16396
rect 37200 16182 37228 16390
rect 37188 16176 37240 16182
rect 37188 16118 37240 16124
rect 37292 16114 37320 17206
rect 37568 16250 37596 18294
rect 37660 17882 37688 19314
rect 37648 17876 37700 17882
rect 37648 17818 37700 17824
rect 37648 17536 37700 17542
rect 37648 17478 37700 17484
rect 37660 17202 37688 17478
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37556 16244 37608 16250
rect 37556 16186 37608 16192
rect 37280 16108 37332 16114
rect 37280 16050 37332 16056
rect 37648 16108 37700 16114
rect 37648 16050 37700 16056
rect 36912 15564 36964 15570
rect 36912 15506 36964 15512
rect 36636 15156 36688 15162
rect 36636 15098 36688 15104
rect 36924 15094 36952 15506
rect 35900 15088 35952 15094
rect 35900 15030 35952 15036
rect 36912 15088 36964 15094
rect 36912 15030 36964 15036
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 34888 15020 34940 15026
rect 34888 14962 34940 14968
rect 35532 15020 35584 15026
rect 35532 14962 35584 14968
rect 32956 14612 33008 14618
rect 32956 14554 33008 14560
rect 33060 14414 33088 14962
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 35544 14618 35572 14962
rect 35532 14612 35584 14618
rect 35532 14554 35584 14560
rect 35912 14482 35940 15030
rect 37292 14618 37320 16050
rect 37660 15502 37688 16050
rect 38292 15904 38344 15910
rect 38292 15846 38344 15852
rect 37648 15496 37700 15502
rect 37648 15438 37700 15444
rect 38108 15428 38160 15434
rect 38108 15370 38160 15376
rect 37648 15360 37700 15366
rect 37648 15302 37700 15308
rect 37660 15026 37688 15302
rect 38120 15162 38148 15370
rect 38108 15156 38160 15162
rect 38108 15098 38160 15104
rect 38304 15026 38332 15846
rect 37648 15020 37700 15026
rect 37648 14962 37700 14968
rect 38292 15020 38344 15026
rect 38292 14962 38344 14968
rect 37464 14816 37516 14822
rect 37464 14758 37516 14764
rect 37280 14612 37332 14618
rect 37280 14554 37332 14560
rect 35900 14476 35952 14482
rect 35900 14418 35952 14424
rect 37476 14414 37504 14758
rect 33048 14408 33100 14414
rect 33048 14350 33100 14356
rect 35440 14408 35492 14414
rect 35440 14350 35492 14356
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 35452 14074 35480 14350
rect 35440 14068 35492 14074
rect 35440 14010 35492 14016
rect 38108 13932 38160 13938
rect 38108 13874 38160 13880
rect 35808 13864 35860 13870
rect 35808 13806 35860 13812
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35820 13394 35848 13806
rect 32772 13388 32824 13394
rect 32772 13330 32824 13336
rect 35808 13388 35860 13394
rect 35808 13330 35860 13336
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 29920 8968 29972 8974
rect 29920 8910 29972 8916
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 38120 2650 38148 13874
rect 38198 8936 38254 8945
rect 38198 8871 38254 8880
rect 38212 8838 38240 8871
rect 38200 8832 38252 8838
rect 38200 8774 38252 8780
rect 29644 2644 29696 2650
rect 29644 2586 29696 2592
rect 38108 2644 38160 2650
rect 38108 2586 38160 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 29000 2440 29052 2446
rect 29000 2382 29052 2388
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 32 800 60 2382
rect 9692 800 9720 2382
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 29012 800 29040 2382
rect 38672 800 38700 2382
rect 18 200 74 800
rect 9678 200 9734 800
rect 19338 200 19394 800
rect 28998 200 29054 800
rect 38658 200 38714 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 1766 30640 1822 30696
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 20258 24148 20260 24168
rect 20260 24148 20312 24168
rect 20312 24148 20314 24168
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 20258 24112 20314 24148
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20810 23024 20866 23080
rect 21914 23060 21916 23080
rect 21916 23060 21968 23080
rect 21968 23060 21970 23080
rect 21914 23024 21970 23060
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 1766 20440 1822 20496
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 1766 10240 1822 10296
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 28906 24112 28962 24168
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 22190 14456 22246 14512
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 28538 15444 28540 15464
rect 28540 15444 28592 15464
rect 28592 15444 28594 15464
rect 28538 15408 28594 15444
rect 28906 15408 28962 15464
rect 27986 14456 28042 14512
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 38290 29280 38346 29336
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34518 19216 34574 19272
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38198 8880 38254 8936
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 200 30698 800 30728
rect 1761 30698 1827 30701
rect 200 30696 1827 30698
rect 200 30640 1766 30696
rect 1822 30640 1827 30696
rect 200 30638 1827 30640
rect 200 30608 800 30638
rect 1761 30635 1827 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 38285 29338 38351 29341
rect 39200 29338 39800 29368
rect 38285 29336 39800 29338
rect 38285 29280 38290 29336
rect 38346 29280 39800 29336
rect 38285 29278 39800 29280
rect 38285 29275 38351 29278
rect 39200 29248 39800 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 20253 24170 20319 24173
rect 28901 24170 28967 24173
rect 20253 24168 28967 24170
rect 20253 24112 20258 24168
rect 20314 24112 28906 24168
rect 28962 24112 28967 24168
rect 20253 24110 28967 24112
rect 20253 24107 20319 24110
rect 28901 24107 28967 24110
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 20805 23082 20871 23085
rect 21909 23082 21975 23085
rect 20805 23080 21975 23082
rect 20805 23024 20810 23080
rect 20866 23024 21914 23080
rect 21970 23024 21975 23080
rect 20805 23022 21975 23024
rect 20805 23019 20871 23022
rect 21909 23019 21975 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 200 20498 800 20528
rect 1761 20498 1827 20501
rect 200 20496 1827 20498
rect 200 20440 1766 20496
rect 1822 20440 1827 20496
rect 200 20438 1827 20440
rect 200 20408 800 20438
rect 1761 20435 1827 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 34513 19274 34579 19277
rect 34513 19272 35910 19274
rect 34513 19216 34518 19272
rect 34574 19216 35910 19272
rect 34513 19214 35910 19216
rect 34513 19211 34579 19214
rect 35850 19138 35910 19214
rect 39200 19138 39800 19168
rect 35850 19078 39800 19138
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 39200 19048 39800 19078
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 28533 15466 28599 15469
rect 28901 15466 28967 15469
rect 28533 15464 28967 15466
rect 28533 15408 28538 15464
rect 28594 15408 28906 15464
rect 28962 15408 28967 15464
rect 28533 15406 28967 15408
rect 28533 15403 28599 15406
rect 28901 15403 28967 15406
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 22185 14514 22251 14517
rect 27981 14514 28047 14517
rect 22185 14512 28047 14514
rect 22185 14456 22190 14512
rect 22246 14456 27986 14512
rect 28042 14456 28047 14512
rect 22185 14454 28047 14456
rect 22185 14451 22251 14454
rect 27981 14451 28047 14454
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 200 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1761 10298 1827 10301
rect 200 10296 1827 10298
rect 200 10240 1766 10296
rect 1822 10240 1827 10296
rect 200 10238 1827 10240
rect 200 10208 800 10238
rect 1761 10235 1827 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 38193 8938 38259 8941
rect 39200 8938 39800 8968
rect 38193 8936 39800 8938
rect 38193 8880 38198 8936
rect 38254 8880 39800 8936
rect 38193 8878 39800 8880
rect 38193 8875 38259 8878
rect 39200 8848 39800 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_1 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 20884 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1667941163
transform 1 0 22816 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1667941163
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1667941163
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1667941163
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1667941163
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1667941163
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_85 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 8924 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1667941163
transform 1 0 9660 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1667941163
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1667941163
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1667941163
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1667941163
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1667941163
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1667941163
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1667941163
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1667941163
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1667941163
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1667941163
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1667941163
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1667941163
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_203
timestamp 1667941163
transform 1 0 19780 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_215
timestamp 1667941163
transform 1 0 20884 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1667941163
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1667941163
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1667941163
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1667941163
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1667941163
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1667941163
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1667941163
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1667941163
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1667941163
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1667941163
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1667941163
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_314
timestamp 1667941163
transform 1 0 29992 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_326
timestamp 1667941163
transform 1 0 31096 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_334
timestamp 1667941163
transform 1 0 31832 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1667941163
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1667941163
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1667941163
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_365
timestamp 1667941163
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_377
timestamp 1667941163
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_389
timestamp 1667941163
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_393
timestamp 1667941163
transform 1 0 37260 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_401
timestamp 1667941163
transform 1 0 37996 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1667941163
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1667941163
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1667941163
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1667941163
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1667941163
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1667941163
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1667941163
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1667941163
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1667941163
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1667941163
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1667941163
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1667941163
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1667941163
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1667941163
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1667941163
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1667941163
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1667941163
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1667941163
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1667941163
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1667941163
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1667941163
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1667941163
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1667941163
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1667941163
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1667941163
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1667941163
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1667941163
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1667941163
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1667941163
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1667941163
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1667941163
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1667941163
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1667941163
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1667941163
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1667941163
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1667941163
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1667941163
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_361
timestamp 1667941163
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_373
timestamp 1667941163
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_385
timestamp 1667941163
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1667941163
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1667941163
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1667941163
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1667941163
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1667941163
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1667941163
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1667941163
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1667941163
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1667941163
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1667941163
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1667941163
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1667941163
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1667941163
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1667941163
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1667941163
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1667941163
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1667941163
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1667941163
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1667941163
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1667941163
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1667941163
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1667941163
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1667941163
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1667941163
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1667941163
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1667941163
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1667941163
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1667941163
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1667941163
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1667941163
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1667941163
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1667941163
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1667941163
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1667941163
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1667941163
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1667941163
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1667941163
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1667941163
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1667941163
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1667941163
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1667941163
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1667941163
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1667941163
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1667941163
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1667941163
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1667941163
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1667941163
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1667941163
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1667941163
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1667941163
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1667941163
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1667941163
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1667941163
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1667941163
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1667941163
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1667941163
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1667941163
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1667941163
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1667941163
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1667941163
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1667941163
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1667941163
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1667941163
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1667941163
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1667941163
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1667941163
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1667941163
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1667941163
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1667941163
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1667941163
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1667941163
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1667941163
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1667941163
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1667941163
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1667941163
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1667941163
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1667941163
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1667941163
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1667941163
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1667941163
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1667941163
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1667941163
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1667941163
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1667941163
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1667941163
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1667941163
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1667941163
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1667941163
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1667941163
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1667941163
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1667941163
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1667941163
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1667941163
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1667941163
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1667941163
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1667941163
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1667941163
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1667941163
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1667941163
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1667941163
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1667941163
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1667941163
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1667941163
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1667941163
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1667941163
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1667941163
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1667941163
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1667941163
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1667941163
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1667941163
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1667941163
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1667941163
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1667941163
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1667941163
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1667941163
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1667941163
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1667941163
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1667941163
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1667941163
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1667941163
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1667941163
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1667941163
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1667941163
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1667941163
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1667941163
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1667941163
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1667941163
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1667941163
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1667941163
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1667941163
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1667941163
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1667941163
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1667941163
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1667941163
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1667941163
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1667941163
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1667941163
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1667941163
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1667941163
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1667941163
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1667941163
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1667941163
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1667941163
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1667941163
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1667941163
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1667941163
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1667941163
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1667941163
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1667941163
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1667941163
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1667941163
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1667941163
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1667941163
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1667941163
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1667941163
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1667941163
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1667941163
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1667941163
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1667941163
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1667941163
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1667941163
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1667941163
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1667941163
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1667941163
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1667941163
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1667941163
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1667941163
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1667941163
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1667941163
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1667941163
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1667941163
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1667941163
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1667941163
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1667941163
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1667941163
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1667941163
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1667941163
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1667941163
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1667941163
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1667941163
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1667941163
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1667941163
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1667941163
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1667941163
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1667941163
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1667941163
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1667941163
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1667941163
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1667941163
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1667941163
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1667941163
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1667941163
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1667941163
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1667941163
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1667941163
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1667941163
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1667941163
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1667941163
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1667941163
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1667941163
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1667941163
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1667941163
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1667941163
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1667941163
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1667941163
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1667941163
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1667941163
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1667941163
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1667941163
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1667941163
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1667941163
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1667941163
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1667941163
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1667941163
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1667941163
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1667941163
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1667941163
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1667941163
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1667941163
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1667941163
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1667941163
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1667941163
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1667941163
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1667941163
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1667941163
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1667941163
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1667941163
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1667941163
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1667941163
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1667941163
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1667941163
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1667941163
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1667941163
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1667941163
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1667941163
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1667941163
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1667941163
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1667941163
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1667941163
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1667941163
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1667941163
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1667941163
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1667941163
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1667941163
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1667941163
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1667941163
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1667941163
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1667941163
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1667941163
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1667941163
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1667941163
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1667941163
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1667941163
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1667941163
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1667941163
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1667941163
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1667941163
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1667941163
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1667941163
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1667941163
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1667941163
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1667941163
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1667941163
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1667941163
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1667941163
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1667941163
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1667941163
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1667941163
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1667941163
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1667941163
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1667941163
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1667941163
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1667941163
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1667941163
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1667941163
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1667941163
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1667941163
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1667941163
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1667941163
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1667941163
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1667941163
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1667941163
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1667941163
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1667941163
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1667941163
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1667941163
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1667941163
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1667941163
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1667941163
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1667941163
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1667941163
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1667941163
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1667941163
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1667941163
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1667941163
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1667941163
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1667941163
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1667941163
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1667941163
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1667941163
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1667941163
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1667941163
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1667941163
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1667941163
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1667941163
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1667941163
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1667941163
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1667941163
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1667941163
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1667941163
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1667941163
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1667941163
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1667941163
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1667941163
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1667941163
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1667941163
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1667941163
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1667941163
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1667941163
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1667941163
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1667941163
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1667941163
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1667941163
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1667941163
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1667941163
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1667941163
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1667941163
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1667941163
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1667941163
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1667941163
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1667941163
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1667941163
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1667941163
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1667941163
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1667941163
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1667941163
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1667941163
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1667941163
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1667941163
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1667941163
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1667941163
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1667941163
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1667941163
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1667941163
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1667941163
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1667941163
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1667941163
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1667941163
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1667941163
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1667941163
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1667941163
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1667941163
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1667941163
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1667941163
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1667941163
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1667941163
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1667941163
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1667941163
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1667941163
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1667941163
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1667941163
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1667941163
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1667941163
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1667941163
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1667941163
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1667941163
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1667941163
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1667941163
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1667941163
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1667941163
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1667941163
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1667941163
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1667941163
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1667941163
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1667941163
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1667941163
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1667941163
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1667941163
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1667941163
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1667941163
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1667941163
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1667941163
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1667941163
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1667941163
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1667941163
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1667941163
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1667941163
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1667941163
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1667941163
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1667941163
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1667941163
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1667941163
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1667941163
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1667941163
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1667941163
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1667941163
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1667941163
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1667941163
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1667941163
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1667941163
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1667941163
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1667941163
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1667941163
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1667941163
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1667941163
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1667941163
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1667941163
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1667941163
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1667941163
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1667941163
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1667941163
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1667941163
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1667941163
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1667941163
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1667941163
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1667941163
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1667941163
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1667941163
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1667941163
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1667941163
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1667941163
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1667941163
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1667941163
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1667941163
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1667941163
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1667941163
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1667941163
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1667941163
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1667941163
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1667941163
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1667941163
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1667941163
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1667941163
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1667941163
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1667941163
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1667941163
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1667941163
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1667941163
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1667941163
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1667941163
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1667941163
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1667941163
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1667941163
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1667941163
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1667941163
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1667941163
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1667941163
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1667941163
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1667941163
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1667941163
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1667941163
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1667941163
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1667941163
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1667941163
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1667941163
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1667941163
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1667941163
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1667941163
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1667941163
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1667941163
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1667941163
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1667941163
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1667941163
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1667941163
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1667941163
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1667941163
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1667941163
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1667941163
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1667941163
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1667941163
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1667941163
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1667941163
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1667941163
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1667941163
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1667941163
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1667941163
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1667941163
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1667941163
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1667941163
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1667941163
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_405
timestamp 1667941163
transform 1 0 38364 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1667941163
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1667941163
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1667941163
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1667941163
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1667941163
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1667941163
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1667941163
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1667941163
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1667941163
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1667941163
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1667941163
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1667941163
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1667941163
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1667941163
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1667941163
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1667941163
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1667941163
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1667941163
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1667941163
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1667941163
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1667941163
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1667941163
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1667941163
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1667941163
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1667941163
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1667941163
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1667941163
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1667941163
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1667941163
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1667941163
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1667941163
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1667941163
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1667941163
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1667941163
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1667941163
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1667941163
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1667941163
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1667941163
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1667941163
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1667941163
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1667941163
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1667941163
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1667941163
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1667941163
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1667941163
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1667941163
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1667941163
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1667941163
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1667941163
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1667941163
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1667941163
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1667941163
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1667941163
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1667941163
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1667941163
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1667941163
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1667941163
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1667941163
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1667941163
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1667941163
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1667941163
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1667941163
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1667941163
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1667941163
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1667941163
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1667941163
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1667941163
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1667941163
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1667941163
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1667941163
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1667941163
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1667941163
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1667941163
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1667941163
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1667941163
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1667941163
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1667941163
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1667941163
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1667941163
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1667941163
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1667941163
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1667941163
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1667941163
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1667941163
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1667941163
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1667941163
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1667941163
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1667941163
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_8
timestamp 1667941163
transform 1 0 1840 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_20
timestamp 1667941163
transform 1 0 2944 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_32
timestamp 1667941163
transform 1 0 4048 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_44
timestamp 1667941163
transform 1 0 5152 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1667941163
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1667941163
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1667941163
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1667941163
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1667941163
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1667941163
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1667941163
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1667941163
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1667941163
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1667941163
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1667941163
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1667941163
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1667941163
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1667941163
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1667941163
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1667941163
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1667941163
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1667941163
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1667941163
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1667941163
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1667941163
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1667941163
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1667941163
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1667941163
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1667941163
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1667941163
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1667941163
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1667941163
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1667941163
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1667941163
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1667941163
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1667941163
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1667941163
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1667941163
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1667941163
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1667941163
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1667941163
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1667941163
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1667941163
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1667941163
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1667941163
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1667941163
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1667941163
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1667941163
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1667941163
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1667941163
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1667941163
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1667941163
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1667941163
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1667941163
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1667941163
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1667941163
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1667941163
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1667941163
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1667941163
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1667941163
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1667941163
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1667941163
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1667941163
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1667941163
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1667941163
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1667941163
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1667941163
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1667941163
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1667941163
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1667941163
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1667941163
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1667941163
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1667941163
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1667941163
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1667941163
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1667941163
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1667941163
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1667941163
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1667941163
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1667941163
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1667941163
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1667941163
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1667941163
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1667941163
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1667941163
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1667941163
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1667941163
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1667941163
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1667941163
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1667941163
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1667941163
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1667941163
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1667941163
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1667941163
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1667941163
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1667941163
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1667941163
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1667941163
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1667941163
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1667941163
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1667941163
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1667941163
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1667941163
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1667941163
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1667941163
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1667941163
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_205
timestamp 1667941163
transform 1 0 19964 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1667941163
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1667941163
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1667941163
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_237
timestamp 1667941163
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_250
timestamp 1667941163
transform 1 0 24104 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_262
timestamp 1667941163
transform 1 0 25208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_274
timestamp 1667941163
transform 1 0 26312 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1667941163
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1667941163
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1667941163
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1667941163
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1667941163
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1667941163
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1667941163
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1667941163
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1667941163
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1667941163
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1667941163
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1667941163
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1667941163
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1667941163
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1667941163
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1667941163
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1667941163
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1667941163
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1667941163
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1667941163
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1667941163
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1667941163
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1667941163
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1667941163
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1667941163
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1667941163
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1667941163
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1667941163
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1667941163
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1667941163
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1667941163
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1667941163
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1667941163
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1667941163
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1667941163
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1667941163
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1667941163
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_205
timestamp 1667941163
transform 1 0 19964 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_216
timestamp 1667941163
transform 1 0 20976 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_223
timestamp 1667941163
transform 1 0 21620 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_234
timestamp 1667941163
transform 1 0 22632 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1667941163
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1667941163
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1667941163
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_265
timestamp 1667941163
transform 1 0 25484 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_269
timestamp 1667941163
transform 1 0 25852 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_277
timestamp 1667941163
transform 1 0 26588 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_283
timestamp 1667941163
transform 1 0 27140 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_287
timestamp 1667941163
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 1667941163
transform 1 0 28612 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1667941163
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1667941163
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1667941163
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1667941163
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1667941163
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1667941163
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1667941163
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1667941163
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1667941163
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1667941163
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_401
timestamp 1667941163
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1667941163
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1667941163
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1667941163
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1667941163
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1667941163
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1667941163
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1667941163
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1667941163
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1667941163
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1667941163
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1667941163
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1667941163
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1667941163
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1667941163
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1667941163
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1667941163
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1667941163
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1667941163
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1667941163
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1667941163
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1667941163
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_205
timestamp 1667941163
transform 1 0 19964 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_212
timestamp 1667941163
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_225
timestamp 1667941163
transform 1 0 21804 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_229
timestamp 1667941163
transform 1 0 22172 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_233
timestamp 1667941163
transform 1 0 22540 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1667941163
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_245
timestamp 1667941163
transform 1 0 23644 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_251
timestamp 1667941163
transform 1 0 24196 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_258
timestamp 1667941163
transform 1 0 24840 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_269
timestamp 1667941163
transform 1 0 25852 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1667941163
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_281
timestamp 1667941163
transform 1 0 26956 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_290
timestamp 1667941163
transform 1 0 27784 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_297
timestamp 1667941163
transform 1 0 28428 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_309
timestamp 1667941163
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_321
timestamp 1667941163
transform 1 0 30636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_333
timestamp 1667941163
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1667941163
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1667941163
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1667941163
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1667941163
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1667941163
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1667941163
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1667941163
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1667941163
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1667941163
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1667941163
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1667941163
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1667941163
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1667941163
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1667941163
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1667941163
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1667941163
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1667941163
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1667941163
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1667941163
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1667941163
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1667941163
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1667941163
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1667941163
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1667941163
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1667941163
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1667941163
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1667941163
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1667941163
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1667941163
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_197
timestamp 1667941163
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1667941163
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_213
timestamp 1667941163
transform 1 0 20700 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_217
timestamp 1667941163
transform 1 0 21068 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_221
timestamp 1667941163
transform 1 0 21436 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_229
timestamp 1667941163
transform 1 0 22172 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_239
timestamp 1667941163
transform 1 0 23092 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_20_249
timestamp 1667941163
transform 1 0 24012 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_253
timestamp 1667941163
transform 1 0 24380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_262
timestamp 1667941163
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_274
timestamp 1667941163
transform 1 0 26312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_282
timestamp 1667941163
transform 1 0 27048 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_293
timestamp 1667941163
transform 1 0 28060 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_297
timestamp 1667941163
transform 1 0 28428 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1667941163
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_309
timestamp 1667941163
transform 1 0 29532 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_316
timestamp 1667941163
transform 1 0 30176 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_328
timestamp 1667941163
transform 1 0 31280 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_340
timestamp 1667941163
transform 1 0 32384 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_352
timestamp 1667941163
transform 1 0 33488 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1667941163
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1667941163
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1667941163
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1667941163
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1667941163
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1667941163
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1667941163
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1667941163
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1667941163
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1667941163
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1667941163
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1667941163
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1667941163
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1667941163
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1667941163
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1667941163
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1667941163
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1667941163
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1667941163
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1667941163
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1667941163
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1667941163
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1667941163
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_181
timestamp 1667941163
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_189
timestamp 1667941163
transform 1 0 18492 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_198
timestamp 1667941163
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_211
timestamp 1667941163
transform 1 0 20516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_219
timestamp 1667941163
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1667941163
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_225
timestamp 1667941163
transform 1 0 21804 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_238
timestamp 1667941163
transform 1 0 23000 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_21_250
timestamp 1667941163
transform 1 0 24104 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_258
timestamp 1667941163
transform 1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_269
timestamp 1667941163
transform 1 0 25852 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_277
timestamp 1667941163
transform 1 0 26588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1667941163
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_21_294
timestamp 1667941163
transform 1 0 28152 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_300
timestamp 1667941163
transform 1 0 28704 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1667941163
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1667941163
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1667941163
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1667941163
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1667941163
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1667941163
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_373
timestamp 1667941163
transform 1 0 35420 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_382
timestamp 1667941163
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1667941163
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1667941163
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1667941163
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1667941163
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1667941163
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1667941163
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1667941163
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1667941163
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1667941163
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1667941163
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1667941163
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1667941163
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1667941163
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1667941163
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1667941163
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1667941163
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1667941163
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1667941163
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1667941163
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1667941163
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1667941163
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1667941163
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1667941163
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1667941163
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1667941163
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_215
timestamp 1667941163
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_227
timestamp 1667941163
transform 1 0 21988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_239
timestamp 1667941163
transform 1 0 23092 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_250
timestamp 1667941163
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1667941163
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_275
timestamp 1667941163
transform 1 0 26404 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_283
timestamp 1667941163
transform 1 0 27140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_291
timestamp 1667941163
transform 1 0 27876 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_300
timestamp 1667941163
transform 1 0 28704 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_22_309
timestamp 1667941163
transform 1 0 29532 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_313
timestamp 1667941163
transform 1 0 29900 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_317
timestamp 1667941163
transform 1 0 30268 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_325
timestamp 1667941163
transform 1 0 31004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_343
timestamp 1667941163
transform 1 0 32660 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_350
timestamp 1667941163
transform 1 0 33304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1667941163
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_22_365
timestamp 1667941163
transform 1 0 34684 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_374
timestamp 1667941163
transform 1 0 35512 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_394
timestamp 1667941163
transform 1 0 37352 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1667941163
transform 1 0 38456 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1667941163
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1667941163
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1667941163
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1667941163
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1667941163
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1667941163
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1667941163
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1667941163
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1667941163
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1667941163
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1667941163
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1667941163
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1667941163
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1667941163
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1667941163
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1667941163
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1667941163
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1667941163
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1667941163
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1667941163
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1667941163
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_205
timestamp 1667941163
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1667941163
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1667941163
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_244
timestamp 1667941163
transform 1 0 23552 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_264
timestamp 1667941163
transform 1 0 25392 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_271
timestamp 1667941163
transform 1 0 26036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_278
timestamp 1667941163
transform 1 0 26680 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_281
timestamp 1667941163
transform 1 0 26956 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_289
timestamp 1667941163
transform 1 0 27692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_298
timestamp 1667941163
transform 1 0 28520 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_305
timestamp 1667941163
transform 1 0 29164 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_313
timestamp 1667941163
transform 1 0 29900 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1667941163
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_337
timestamp 1667941163
transform 1 0 32108 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_343
timestamp 1667941163
transform 1 0 32660 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_349
timestamp 1667941163
transform 1 0 33212 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_369
timestamp 1667941163
transform 1 0 35052 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_23_389
timestamp 1667941163
transform 1 0 36892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1667941163
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_398
timestamp 1667941163
transform 1 0 37720 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1667941163
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1667941163
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1667941163
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1667941163
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1667941163
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1667941163
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1667941163
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1667941163
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1667941163
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1667941163
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1667941163
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1667941163
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1667941163
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1667941163
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1667941163
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1667941163
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1667941163
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1667941163
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1667941163
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1667941163
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1667941163
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1667941163
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1667941163
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_212
timestamp 1667941163
transform 1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_220
timestamp 1667941163
transform 1 0 21344 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_24_231
timestamp 1667941163
transform 1 0 22356 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_240
timestamp 1667941163
transform 1 0 23184 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_247
timestamp 1667941163
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1667941163
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1667941163
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1667941163
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_277
timestamp 1667941163
transform 1 0 26588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_282
timestamp 1667941163
transform 1 0 27048 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_290
timestamp 1667941163
transform 1 0 27784 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_296
timestamp 1667941163
transform 1 0 28336 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_305
timestamp 1667941163
transform 1 0 29164 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_24_309
timestamp 1667941163
transform 1 0 29532 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_318
timestamp 1667941163
transform 1 0 30360 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_325
timestamp 1667941163
transform 1 0 31004 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_334
timestamp 1667941163
transform 1 0 31832 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_342
timestamp 1667941163
transform 1 0 32568 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_351
timestamp 1667941163
transform 1 0 33396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1667941163
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_365
timestamp 1667941163
transform 1 0 34684 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_370
timestamp 1667941163
transform 1 0 35144 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_378
timestamp 1667941163
transform 1 0 35880 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_385
timestamp 1667941163
transform 1 0 36524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_405
timestamp 1667941163
transform 1 0 38364 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1667941163
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1667941163
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1667941163
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1667941163
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1667941163
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1667941163
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1667941163
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1667941163
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1667941163
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1667941163
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1667941163
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1667941163
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1667941163
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1667941163
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1667941163
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1667941163
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1667941163
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1667941163
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1667941163
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1667941163
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1667941163
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_25_207
timestamp 1667941163
transform 1 0 20148 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1667941163
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_225
timestamp 1667941163
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_234
timestamp 1667941163
transform 1 0 22632 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_238
timestamp 1667941163
transform 1 0 23000 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_244
timestamp 1667941163
transform 1 0 23552 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_261
timestamp 1667941163
transform 1 0 25116 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_272
timestamp 1667941163
transform 1 0 26128 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1667941163
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_289
timestamp 1667941163
transform 1 0 27692 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_296
timestamp 1667941163
transform 1 0 28336 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_316
timestamp 1667941163
transform 1 0 30176 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_323
timestamp 1667941163
transform 1 0 30820 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_334
timestamp 1667941163
transform 1 0 31832 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_337
timestamp 1667941163
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_350
timestamp 1667941163
transform 1 0 33304 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_360
timestamp 1667941163
transform 1 0 34224 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_372
timestamp 1667941163
transform 1 0 35328 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_378
timestamp 1667941163
transform 1 0 35880 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_382
timestamp 1667941163
transform 1 0 36248 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_390
timestamp 1667941163
transform 1 0 36984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_393
timestamp 1667941163
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_400
timestamp 1667941163
transform 1 0 37904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_406
timestamp 1667941163
transform 1 0 38456 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1667941163
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1667941163
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1667941163
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1667941163
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1667941163
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1667941163
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1667941163
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1667941163
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1667941163
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1667941163
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1667941163
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1667941163
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1667941163
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1667941163
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1667941163
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1667941163
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1667941163
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1667941163
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1667941163
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1667941163
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1667941163
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1667941163
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_205
timestamp 1667941163
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_26_217
timestamp 1667941163
transform 1 0 21068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_225
timestamp 1667941163
transform 1 0 21804 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_236
timestamp 1667941163
transform 1 0 22816 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_247
timestamp 1667941163
transform 1 0 23828 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1667941163
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1667941163
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_268
timestamp 1667941163
transform 1 0 25760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_292
timestamp 1667941163
transform 1 0 27968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_299
timestamp 1667941163
transform 1 0 28612 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_306
timestamp 1667941163
transform 1 0 29256 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_309
timestamp 1667941163
transform 1 0 29532 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_315
timestamp 1667941163
transform 1 0 30084 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_332
timestamp 1667941163
transform 1 0 31648 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_352
timestamp 1667941163
transform 1 0 33488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1667941163
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_365
timestamp 1667941163
transform 1 0 34684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_383
timestamp 1667941163
transform 1 0 36340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_405
timestamp 1667941163
transform 1 0 38364 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1667941163
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1667941163
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1667941163
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1667941163
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1667941163
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1667941163
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1667941163
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1667941163
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1667941163
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1667941163
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1667941163
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1667941163
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1667941163
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1667941163
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1667941163
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1667941163
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1667941163
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1667941163
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1667941163
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1667941163
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_193
timestamp 1667941163
transform 1 0 18860 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1667941163
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_216
timestamp 1667941163
transform 1 0 20976 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_27_225
timestamp 1667941163
transform 1 0 21804 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_233
timestamp 1667941163
transform 1 0 22540 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_238
timestamp 1667941163
transform 1 0 23000 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_262
timestamp 1667941163
transform 1 0 25208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_270
timestamp 1667941163
transform 1 0 25944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_278
timestamp 1667941163
transform 1 0 26680 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_281
timestamp 1667941163
transform 1 0 26956 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_287
timestamp 1667941163
transform 1 0 27508 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_295
timestamp 1667941163
transform 1 0 28244 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_312
timestamp 1667941163
transform 1 0 29808 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1667941163
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_337
timestamp 1667941163
transform 1 0 32108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_346
timestamp 1667941163
transform 1 0 32936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_350
timestamp 1667941163
transform 1 0 33304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_367
timestamp 1667941163
transform 1 0 34868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_374
timestamp 1667941163
transform 1 0 35512 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_382
timestamp 1667941163
transform 1 0 36248 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1667941163
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_393
timestamp 1667941163
transform 1 0 37260 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_398
timestamp 1667941163
transform 1 0 37720 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_406
timestamp 1667941163
transform 1 0 38456 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1667941163
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1667941163
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1667941163
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1667941163
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1667941163
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1667941163
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1667941163
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1667941163
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1667941163
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1667941163
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1667941163
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1667941163
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1667941163
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1667941163
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1667941163
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1667941163
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1667941163
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1667941163
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1667941163
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1667941163
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1667941163
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1667941163
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_211
timestamp 1667941163
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_219
timestamp 1667941163
transform 1 0 21252 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_227
timestamp 1667941163
transform 1 0 21988 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_235
timestamp 1667941163
transform 1 0 22724 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_244
timestamp 1667941163
transform 1 0 23552 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_253
timestamp 1667941163
transform 1 0 24380 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_264
timestamp 1667941163
transform 1 0 25392 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_273
timestamp 1667941163
transform 1 0 26220 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_282
timestamp 1667941163
transform 1 0 27048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_291
timestamp 1667941163
transform 1 0 27876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_299
timestamp 1667941163
transform 1 0 28612 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_305
timestamp 1667941163
transform 1 0 29164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_309
timestamp 1667941163
transform 1 0 29532 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_314
timestamp 1667941163
transform 1 0 29992 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_323
timestamp 1667941163
transform 1 0 30820 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_347
timestamp 1667941163
transform 1 0 33028 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_356
timestamp 1667941163
transform 1 0 33856 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_28_365
timestamp 1667941163
transform 1 0 34684 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_28_378
timestamp 1667941163
transform 1 0 35880 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_384
timestamp 1667941163
transform 1 0 36432 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_390
timestamp 1667941163
transform 1 0 36984 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_399
timestamp 1667941163
transform 1 0 37812 0 1 17408
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1667941163
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1667941163
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1667941163
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1667941163
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1667941163
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1667941163
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1667941163
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1667941163
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1667941163
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1667941163
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1667941163
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1667941163
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1667941163
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1667941163
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1667941163
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1667941163
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1667941163
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1667941163
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1667941163
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1667941163
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_193
timestamp 1667941163
transform 1 0 18860 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_201
timestamp 1667941163
transform 1 0 19596 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_208
timestamp 1667941163
transform 1 0 20240 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1667941163
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1667941163
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_225
timestamp 1667941163
transform 1 0 21804 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_235
timestamp 1667941163
transform 1 0 22724 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_241
timestamp 1667941163
transform 1 0 23276 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_262
timestamp 1667941163
transform 1 0 25208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_272
timestamp 1667941163
transform 1 0 26128 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_281
timestamp 1667941163
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_299
timestamp 1667941163
transform 1 0 28612 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_327
timestamp 1667941163
transform 1 0 31188 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1667941163
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_337
timestamp 1667941163
transform 1 0 32108 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_356
timestamp 1667941163
transform 1 0 33856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_370
timestamp 1667941163
transform 1 0 35144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_374
timestamp 1667941163
transform 1 0 35512 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_380
timestamp 1667941163
transform 1 0 36064 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_389
timestamp 1667941163
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_393
timestamp 1667941163
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_400
timestamp 1667941163
transform 1 0 37904 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_406
timestamp 1667941163
transform 1 0 38456 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1667941163
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1667941163
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1667941163
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1667941163
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1667941163
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1667941163
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1667941163
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1667941163
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1667941163
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1667941163
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1667941163
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1667941163
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1667941163
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1667941163
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1667941163
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1667941163
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1667941163
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1667941163
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1667941163
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1667941163
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1667941163
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1667941163
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_217
timestamp 1667941163
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_226
timestamp 1667941163
transform 1 0 21896 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_232
timestamp 1667941163
transform 1 0 22448 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_249
timestamp 1667941163
transform 1 0 24012 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 1667941163
transform 1 0 24380 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_271
timestamp 1667941163
transform 1 0 26036 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_291
timestamp 1667941163
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_30_302
timestamp 1667941163
transform 1 0 28888 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1667941163
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_321
timestamp 1667941163
transform 1 0 30636 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_30_347
timestamp 1667941163
transform 1 0 33028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_354
timestamp 1667941163
transform 1 0 33672 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_361
timestamp 1667941163
transform 1 0 34316 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_365
timestamp 1667941163
transform 1 0 34684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_383
timestamp 1667941163
transform 1 0 36340 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1667941163
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1667941163
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1667941163
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1667941163
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1667941163
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1667941163
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1667941163
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1667941163
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1667941163
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1667941163
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1667941163
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1667941163
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1667941163
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1667941163
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1667941163
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1667941163
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1667941163
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1667941163
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1667941163
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1667941163
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1667941163
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_193
timestamp 1667941163
transform 1 0 18860 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_201
timestamp 1667941163
transform 1 0 19596 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_205
timestamp 1667941163
transform 1 0 19964 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_215
timestamp 1667941163
transform 1 0 20884 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1667941163
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_225
timestamp 1667941163
transform 1 0 21804 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_243
timestamp 1667941163
transform 1 0 23460 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1667941163
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1667941163
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_281
timestamp 1667941163
transform 1 0 26956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_286
timestamp 1667941163
transform 1 0 27416 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_31_300
timestamp 1667941163
transform 1 0 28704 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_309
timestamp 1667941163
transform 1 0 29532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_316
timestamp 1667941163
transform 1 0 30176 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_325
timestamp 1667941163
transform 1 0 31004 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_334
timestamp 1667941163
transform 1 0 31832 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_337
timestamp 1667941163
transform 1 0 32108 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_345
timestamp 1667941163
transform 1 0 32844 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_354
timestamp 1667941163
transform 1 0 33672 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_362
timestamp 1667941163
transform 1 0 34408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_366
timestamp 1667941163
transform 1 0 34776 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1667941163
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_393
timestamp 1667941163
transform 1 0 37260 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_398
timestamp 1667941163
transform 1 0 37720 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_406
timestamp 1667941163
transform 1 0 38456 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1667941163
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1667941163
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1667941163
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1667941163
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1667941163
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1667941163
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1667941163
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1667941163
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1667941163
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1667941163
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1667941163
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1667941163
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1667941163
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1667941163
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1667941163
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1667941163
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1667941163
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1667941163
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1667941163
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1667941163
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1667941163
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1667941163
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_203
timestamp 1667941163
transform 1 0 19780 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_220
timestamp 1667941163
transform 1 0 21344 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_228
timestamp 1667941163
transform 1 0 22080 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_232
timestamp 1667941163
transform 1 0 22448 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_244
timestamp 1667941163
transform 1 0 23552 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1667941163
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_253
timestamp 1667941163
transform 1 0 24380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_257
timestamp 1667941163
transform 1 0 24748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_262
timestamp 1667941163
transform 1 0 25208 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_268
timestamp 1667941163
transform 1 0 25760 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_274
timestamp 1667941163
transform 1 0 26312 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_286
timestamp 1667941163
transform 1 0 27416 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_294
timestamp 1667941163
transform 1 0 28152 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_300
timestamp 1667941163
transform 1 0 28704 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_309
timestamp 1667941163
transform 1 0 29532 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_316
timestamp 1667941163
transform 1 0 30176 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_324
timestamp 1667941163
transform 1 0 30912 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_331
timestamp 1667941163
transform 1 0 31556 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_339
timestamp 1667941163
transform 1 0 32292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1667941163
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1667941163
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_365
timestamp 1667941163
transform 1 0 34684 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_372
timestamp 1667941163
transform 1 0 35328 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_376
timestamp 1667941163
transform 1 0 35696 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_380
timestamp 1667941163
transform 1 0 36064 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_392
timestamp 1667941163
transform 1 0 37168 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_404
timestamp 1667941163
transform 1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1667941163
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1667941163
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1667941163
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1667941163
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1667941163
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1667941163
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1667941163
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1667941163
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1667941163
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1667941163
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1667941163
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1667941163
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1667941163
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1667941163
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1667941163
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1667941163
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1667941163
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1667941163
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1667941163
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1667941163
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_193
timestamp 1667941163
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_207
timestamp 1667941163
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_214
timestamp 1667941163
transform 1 0 20792 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_222
timestamp 1667941163
transform 1 0 21528 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1667941163
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1667941163
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_249
timestamp 1667941163
transform 1 0 24012 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_255
timestamp 1667941163
transform 1 0 24564 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_261
timestamp 1667941163
transform 1 0 25116 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_278
timestamp 1667941163
transform 1 0 26680 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1667941163
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_296
timestamp 1667941163
transform 1 0 28336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_316
timestamp 1667941163
transform 1 0 30176 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1667941163
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1667941163
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_337
timestamp 1667941163
transform 1 0 32108 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_345
timestamp 1667941163
transform 1 0 32844 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_354
timestamp 1667941163
transform 1 0 33672 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_361
timestamp 1667941163
transform 1 0 34316 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_369
timestamp 1667941163
transform 1 0 35052 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_375
timestamp 1667941163
transform 1 0 35604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_382
timestamp 1667941163
transform 1 0 36248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1667941163
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1667941163
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1667941163
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_3
timestamp 1667941163
transform 1 0 1380 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_8
timestamp 1667941163
transform 1 0 1840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1667941163
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1667941163
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1667941163
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1667941163
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1667941163
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1667941163
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1667941163
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1667941163
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1667941163
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1667941163
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1667941163
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1667941163
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1667941163
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1667941163
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1667941163
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1667941163
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1667941163
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1667941163
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1667941163
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1667941163
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1667941163
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_221
timestamp 1667941163
transform 1 0 21436 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_229
timestamp 1667941163
transform 1 0 22172 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1667941163
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_253
timestamp 1667941163
transform 1 0 24380 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1667941163
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1667941163
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_302
timestamp 1667941163
transform 1 0 28888 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_309
timestamp 1667941163
transform 1 0 29532 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_34_333
timestamp 1667941163
transform 1 0 31740 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_341
timestamp 1667941163
transform 1 0 32476 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_359
timestamp 1667941163
transform 1 0 34132 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1667941163
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_365
timestamp 1667941163
transform 1 0 34684 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_383
timestamp 1667941163
transform 1 0 36340 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_395
timestamp 1667941163
transform 1 0 37444 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1667941163
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1667941163
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1667941163
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1667941163
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1667941163
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1667941163
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1667941163
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1667941163
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1667941163
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1667941163
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1667941163
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1667941163
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1667941163
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1667941163
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1667941163
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1667941163
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1667941163
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1667941163
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1667941163
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_181
timestamp 1667941163
transform 1 0 17756 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_189
timestamp 1667941163
transform 1 0 18492 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_194
timestamp 1667941163
transform 1 0 18952 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_202
timestamp 1667941163
transform 1 0 19688 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1667941163
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1667941163
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_225
timestamp 1667941163
transform 1 0 21804 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1667941163
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_250
timestamp 1667941163
transform 1 0 24104 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_262
timestamp 1667941163
transform 1 0 25208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_266
timestamp 1667941163
transform 1 0 25576 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_270
timestamp 1667941163
transform 1 0 25944 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_274
timestamp 1667941163
transform 1 0 26312 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_278
timestamp 1667941163
transform 1 0 26680 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_281
timestamp 1667941163
transform 1 0 26956 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_288
timestamp 1667941163
transform 1 0 27600 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_299
timestamp 1667941163
transform 1 0 28612 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_308
timestamp 1667941163
transform 1 0 29440 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_320
timestamp 1667941163
transform 1 0 30544 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_328
timestamp 1667941163
transform 1 0 31280 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_337
timestamp 1667941163
transform 1 0 32108 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_347
timestamp 1667941163
transform 1 0 33028 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_355
timestamp 1667941163
transform 1 0 33764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_361
timestamp 1667941163
transform 1 0 34316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_367
timestamp 1667941163
transform 1 0 34868 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_387
timestamp 1667941163
transform 1 0 36708 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1667941163
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1667941163
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1667941163
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1667941163
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1667941163
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1667941163
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1667941163
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1667941163
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1667941163
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1667941163
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1667941163
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1667941163
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1667941163
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1667941163
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1667941163
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1667941163
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1667941163
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1667941163
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1667941163
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1667941163
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1667941163
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_177
timestamp 1667941163
transform 1 0 17388 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_184
timestamp 1667941163
transform 1 0 18032 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1667941163
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_197
timestamp 1667941163
transform 1 0 19228 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_205
timestamp 1667941163
transform 1 0 19964 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_212
timestamp 1667941163
transform 1 0 20608 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_220
timestamp 1667941163
transform 1 0 21344 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1667941163
transform 1 0 22632 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_242
timestamp 1667941163
transform 1 0 23368 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_250
timestamp 1667941163
transform 1 0 24104 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_253
timestamp 1667941163
transform 1 0 24380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_260
timestamp 1667941163
transform 1 0 25024 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_266
timestamp 1667941163
transform 1 0 25576 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_272
timestamp 1667941163
transform 1 0 26128 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_282
timestamp 1667941163
transform 1 0 27048 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_294
timestamp 1667941163
transform 1 0 28152 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_299
timestamp 1667941163
transform 1 0 28612 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_306
timestamp 1667941163
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_309
timestamp 1667941163
transform 1 0 29532 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_313
timestamp 1667941163
transform 1 0 29900 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_330
timestamp 1667941163
transform 1 0 31464 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_336
timestamp 1667941163
transform 1 0 32016 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_344
timestamp 1667941163
transform 1 0 32752 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_352
timestamp 1667941163
transform 1 0 33488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_356
timestamp 1667941163
transform 1 0 33856 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_362
timestamp 1667941163
transform 1 0 34408 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_365
timestamp 1667941163
transform 1 0 34684 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_375
timestamp 1667941163
transform 1 0 35604 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_385
timestamp 1667941163
transform 1 0 36524 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_393
timestamp 1667941163
transform 1 0 37260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_397
timestamp 1667941163
transform 1 0 37628 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_405
timestamp 1667941163
transform 1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1667941163
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1667941163
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1667941163
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1667941163
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1667941163
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1667941163
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1667941163
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1667941163
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1667941163
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1667941163
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1667941163
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1667941163
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1667941163
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1667941163
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1667941163
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1667941163
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1667941163
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1667941163
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_169
timestamp 1667941163
transform 1 0 16652 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_177
timestamp 1667941163
transform 1 0 17388 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_185
timestamp 1667941163
transform 1 0 18124 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_197
timestamp 1667941163
transform 1 0 19228 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1667941163
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1667941163
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_225
timestamp 1667941163
transform 1 0 21804 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1667941163
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_246
timestamp 1667941163
transform 1 0 23736 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_268
timestamp 1667941163
transform 1 0 25760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_278
timestamp 1667941163
transform 1 0 26680 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1667941163
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_305
timestamp 1667941163
transform 1 0 29164 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_312
timestamp 1667941163
transform 1 0 29808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_322
timestamp 1667941163
transform 1 0 30728 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1667941163
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1667941163
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_337
timestamp 1667941163
transform 1 0 32108 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_355
timestamp 1667941163
transform 1 0 33764 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_359
timestamp 1667941163
transform 1 0 34132 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_363
timestamp 1667941163
transform 1 0 34500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_383
timestamp 1667941163
transform 1 0 36340 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1667941163
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_393
timestamp 1667941163
transform 1 0 37260 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_37_400
timestamp 1667941163
transform 1 0 37904 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_406
timestamp 1667941163
transform 1 0 38456 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1667941163
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1667941163
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1667941163
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1667941163
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1667941163
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1667941163
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1667941163
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1667941163
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1667941163
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1667941163
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1667941163
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1667941163
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1667941163
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1667941163
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1667941163
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1667941163
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1667941163
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1667941163
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1667941163
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_184
timestamp 1667941163
transform 1 0 18032 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1667941163
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_197
timestamp 1667941163
transform 1 0 19228 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1667941163
transform 1 0 19780 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_211
timestamp 1667941163
transform 1 0 20516 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_216
timestamp 1667941163
transform 1 0 20976 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_227
timestamp 1667941163
transform 1 0 21988 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_233
timestamp 1667941163
transform 1 0 22540 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_250
timestamp 1667941163
transform 1 0 24104 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_253
timestamp 1667941163
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_264
timestamp 1667941163
transform 1 0 25392 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_276
timestamp 1667941163
transform 1 0 26496 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_283
timestamp 1667941163
transform 1 0 27140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_287
timestamp 1667941163
transform 1 0 27508 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1667941163
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_38_309
timestamp 1667941163
transform 1 0 29532 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_331
timestamp 1667941163
transform 1 0 31556 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_340
timestamp 1667941163
transform 1 0 32384 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_352
timestamp 1667941163
transform 1 0 33488 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_38_361
timestamp 1667941163
transform 1 0 34316 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_365
timestamp 1667941163
transform 1 0 34684 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_383
timestamp 1667941163
transform 1 0 36340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_38_405
timestamp 1667941163
transform 1 0 38364 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1667941163
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1667941163
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1667941163
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1667941163
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1667941163
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1667941163
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1667941163
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1667941163
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1667941163
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1667941163
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1667941163
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1667941163
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1667941163
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1667941163
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1667941163
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1667941163
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1667941163
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1667941163
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1667941163
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_187
timestamp 1667941163
transform 1 0 18308 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_195
timestamp 1667941163
transform 1 0 19044 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_39_200
timestamp 1667941163
transform 1 0 19504 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_212
timestamp 1667941163
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_218
timestamp 1667941163
transform 1 0 21160 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_222
timestamp 1667941163
transform 1 0 21528 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_225
timestamp 1667941163
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_236
timestamp 1667941163
transform 1 0 22816 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_262
timestamp 1667941163
transform 1 0 25208 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_275
timestamp 1667941163
transform 1 0 26404 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1667941163
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1667941163
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_293
timestamp 1667941163
transform 1 0 28060 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_301
timestamp 1667941163
transform 1 0 28796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_306
timestamp 1667941163
transform 1 0 29256 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_314
timestamp 1667941163
transform 1 0 29992 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1667941163
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1667941163
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1667941163
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_349
timestamp 1667941163
transform 1 0 33212 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_375
timestamp 1667941163
transform 1 0 35604 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_383
timestamp 1667941163
transform 1 0 36340 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_39_389
timestamp 1667941163
transform 1 0 36892 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_39_393
timestamp 1667941163
transform 1 0 37260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_39_400
timestamp 1667941163
transform 1 0 37904 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_406
timestamp 1667941163
transform 1 0 38456 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1667941163
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1667941163
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1667941163
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1667941163
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1667941163
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1667941163
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1667941163
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1667941163
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1667941163
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1667941163
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1667941163
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1667941163
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1667941163
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1667941163
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1667941163
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1667941163
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1667941163
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_165
timestamp 1667941163
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_171
timestamp 1667941163
transform 1 0 16836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_176
timestamp 1667941163
transform 1 0 17296 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_187
timestamp 1667941163
transform 1 0 18308 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_194
timestamp 1667941163
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_197
timestamp 1667941163
transform 1 0 19228 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_208
timestamp 1667941163
transform 1 0 20240 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_219
timestamp 1667941163
transform 1 0 21252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_231
timestamp 1667941163
transform 1 0 22356 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_242
timestamp 1667941163
transform 1 0 23368 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_250
timestamp 1667941163
transform 1 0 24104 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_253
timestamp 1667941163
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_258
timestamp 1667941163
transform 1 0 24840 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_262
timestamp 1667941163
transform 1 0 25208 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_279
timestamp 1667941163
transform 1 0 26772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_287
timestamp 1667941163
transform 1 0 27508 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_295
timestamp 1667941163
transform 1 0 28244 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1667941163
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_309
timestamp 1667941163
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_316
timestamp 1667941163
transform 1 0 30176 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1667941163
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_332
timestamp 1667941163
transform 1 0 31648 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_352
timestamp 1667941163
transform 1 0 33488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_40_361
timestamp 1667941163
transform 1 0 34316 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_365
timestamp 1667941163
transform 1 0 34684 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_370
timestamp 1667941163
transform 1 0 35144 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_378
timestamp 1667941163
transform 1 0 35880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_397
timestamp 1667941163
transform 1 0 37628 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_405
timestamp 1667941163
transform 1 0 38364 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1667941163
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1667941163
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1667941163
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1667941163
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1667941163
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1667941163
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1667941163
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1667941163
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1667941163
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1667941163
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1667941163
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1667941163
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1667941163
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1667941163
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1667941163
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1667941163
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_161
timestamp 1667941163
transform 1 0 15916 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1667941163
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1667941163
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1667941163
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_186
timestamp 1667941163
transform 1 0 18216 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_196
timestamp 1667941163
transform 1 0 19136 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1667941163
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_225
timestamp 1667941163
transform 1 0 21804 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_232
timestamp 1667941163
transform 1 0 22448 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1667941163
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_259
timestamp 1667941163
transform 1 0 24932 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_266
timestamp 1667941163
transform 1 0 25576 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1667941163
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_281
timestamp 1667941163
transform 1 0 26956 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_299
timestamp 1667941163
transform 1 0 28612 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_319
timestamp 1667941163
transform 1 0 30452 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_326
timestamp 1667941163
transform 1 0 31096 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_41_333
timestamp 1667941163
transform 1 0 31740 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_337
timestamp 1667941163
transform 1 0 32108 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_341
timestamp 1667941163
transform 1 0 32476 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_348
timestamp 1667941163
transform 1 0 33120 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_355
timestamp 1667941163
transform 1 0 33764 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_370
timestamp 1667941163
transform 1 0 35144 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_382
timestamp 1667941163
transform 1 0 36248 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_390
timestamp 1667941163
transform 1 0 36984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_393
timestamp 1667941163
transform 1 0 37260 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_402
timestamp 1667941163
transform 1 0 38088 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_406
timestamp 1667941163
transform 1 0 38456 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1667941163
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1667941163
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1667941163
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1667941163
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1667941163
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1667941163
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1667941163
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1667941163
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1667941163
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1667941163
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1667941163
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1667941163
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1667941163
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1667941163
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1667941163
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1667941163
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1667941163
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_165
timestamp 1667941163
transform 1 0 16284 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_173
timestamp 1667941163
transform 1 0 17020 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_182
timestamp 1667941163
transform 1 0 17848 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_194
timestamp 1667941163
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_197
timestamp 1667941163
transform 1 0 19228 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_219
timestamp 1667941163
transform 1 0 21252 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_230
timestamp 1667941163
transform 1 0 22264 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1667941163
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1667941163
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1667941163
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_267
timestamp 1667941163
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_271
timestamp 1667941163
transform 1 0 26036 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_277
timestamp 1667941163
transform 1 0 26588 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_286
timestamp 1667941163
transform 1 0 27416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_293
timestamp 1667941163
transform 1 0 28060 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_306
timestamp 1667941163
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1667941163
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_313
timestamp 1667941163
transform 1 0 29900 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_330
timestamp 1667941163
transform 1 0 31464 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_352
timestamp 1667941163
transform 1 0 33488 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1667941163
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_365
timestamp 1667941163
transform 1 0 34684 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_383
timestamp 1667941163
transform 1 0 36340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_405
timestamp 1667941163
transform 1 0 38364 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1667941163
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1667941163
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1667941163
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1667941163
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1667941163
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1667941163
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1667941163
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1667941163
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1667941163
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1667941163
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1667941163
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1667941163
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1667941163
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1667941163
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1667941163
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1667941163
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1667941163
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1667941163
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_169
timestamp 1667941163
transform 1 0 16652 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_43_184
timestamp 1667941163
transform 1 0 18032 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_196
timestamp 1667941163
transform 1 0 19136 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_43_207
timestamp 1667941163
transform 1 0 20148 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_219
timestamp 1667941163
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1667941163
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_225
timestamp 1667941163
transform 1 0 21804 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_238
timestamp 1667941163
transform 1 0 23000 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_262
timestamp 1667941163
transform 1 0 25208 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_270
timestamp 1667941163
transform 1 0 25944 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_278
timestamp 1667941163
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1667941163
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_293
timestamp 1667941163
transform 1 0 28060 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_301
timestamp 1667941163
transform 1 0 28796 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_308
timestamp 1667941163
transform 1 0 29440 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_328
timestamp 1667941163
transform 1 0 31280 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_337
timestamp 1667941163
transform 1 0 32108 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_342
timestamp 1667941163
transform 1 0 32568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_362
timestamp 1667941163
transform 1 0 34408 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_371
timestamp 1667941163
transform 1 0 35236 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_379
timestamp 1667941163
transform 1 0 35972 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_383
timestamp 1667941163
transform 1 0 36340 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1667941163
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_393
timestamp 1667941163
transform 1 0 37260 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_400
timestamp 1667941163
transform 1 0 37904 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_406
timestamp 1667941163
transform 1 0 38456 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1667941163
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1667941163
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1667941163
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1667941163
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1667941163
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1667941163
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1667941163
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1667941163
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1667941163
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1667941163
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1667941163
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1667941163
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1667941163
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1667941163
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1667941163
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1667941163
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1667941163
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1667941163
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_177
timestamp 1667941163
transform 1 0 17388 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_181
timestamp 1667941163
transform 1 0 17756 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_185
timestamp 1667941163
transform 1 0 18124 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_193
timestamp 1667941163
transform 1 0 18860 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1667941163
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_209
timestamp 1667941163
transform 1 0 20332 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_217
timestamp 1667941163
transform 1 0 21068 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_222
timestamp 1667941163
transform 1 0 21528 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_234
timestamp 1667941163
transform 1 0 22632 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_44_240
timestamp 1667941163
transform 1 0 23184 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_253
timestamp 1667941163
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_44_277
timestamp 1667941163
transform 1 0 26588 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_288
timestamp 1667941163
transform 1 0 27600 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_295
timestamp 1667941163
transform 1 0 28244 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_301
timestamp 1667941163
transform 1 0 28796 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_44_305
timestamp 1667941163
transform 1 0 29164 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1667941163
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_319
timestamp 1667941163
transform 1 0 30452 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_347
timestamp 1667941163
transform 1 0 33028 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_356
timestamp 1667941163
transform 1 0 33856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_365
timestamp 1667941163
transform 1 0 34684 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_375
timestamp 1667941163
transform 1 0 35604 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_379
timestamp 1667941163
transform 1 0 35972 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_385
timestamp 1667941163
transform 1 0 36524 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_405
timestamp 1667941163
transform 1 0 38364 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1667941163
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1667941163
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1667941163
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1667941163
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1667941163
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1667941163
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1667941163
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1667941163
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1667941163
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1667941163
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1667941163
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1667941163
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1667941163
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1667941163
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1667941163
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1667941163
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1667941163
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1667941163
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1667941163
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1667941163
transform 1 0 17388 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_186
timestamp 1667941163
transform 1 0 18216 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1667941163
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_218
timestamp 1667941163
transform 1 0 21160 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_45_225
timestamp 1667941163
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_45_236
timestamp 1667941163
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_264
timestamp 1667941163
transform 1 0 25392 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1667941163
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_281
timestamp 1667941163
transform 1 0 26956 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_286
timestamp 1667941163
transform 1 0 27416 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_302
timestamp 1667941163
transform 1 0 28888 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_308
timestamp 1667941163
transform 1 0 29440 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_313
timestamp 1667941163
transform 1 0 29900 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_321
timestamp 1667941163
transform 1 0 30636 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_329
timestamp 1667941163
transform 1 0 31372 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_334
timestamp 1667941163
transform 1 0 31832 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_337
timestamp 1667941163
transform 1 0 32108 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_45_346
timestamp 1667941163
transform 1 0 32936 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_357
timestamp 1667941163
transform 1 0 33948 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_377
timestamp 1667941163
transform 1 0 35788 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_388
timestamp 1667941163
transform 1 0 36800 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_393
timestamp 1667941163
transform 1 0 37260 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_400
timestamp 1667941163
transform 1 0 37904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_406
timestamp 1667941163
transform 1 0 38456 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1667941163
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1667941163
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1667941163
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1667941163
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1667941163
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1667941163
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1667941163
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1667941163
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1667941163
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1667941163
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1667941163
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1667941163
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1667941163
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1667941163
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1667941163
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1667941163
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1667941163
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_172
timestamp 1667941163
transform 1 0 16928 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1667941163
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_191
timestamp 1667941163
transform 1 0 18676 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1667941163
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1667941163
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1667941163
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_221
timestamp 1667941163
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_240
timestamp 1667941163
transform 1 0 23184 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_247
timestamp 1667941163
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1667941163
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_253
timestamp 1667941163
transform 1 0 24380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_258
timestamp 1667941163
transform 1 0 24840 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_266
timestamp 1667941163
transform 1 0 25576 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_271
timestamp 1667941163
transform 1 0 26036 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_275
timestamp 1667941163
transform 1 0 26404 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_283
timestamp 1667941163
transform 1 0 27140 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_296
timestamp 1667941163
transform 1 0 28336 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_302
timestamp 1667941163
transform 1 0 28888 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_46_306
timestamp 1667941163
transform 1 0 29256 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_309
timestamp 1667941163
transform 1 0 29532 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_320
timestamp 1667941163
transform 1 0 30544 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_326
timestamp 1667941163
transform 1 0 31096 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_343
timestamp 1667941163
transform 1 0 32660 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_353
timestamp 1667941163
transform 1 0 33580 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1667941163
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_365
timestamp 1667941163
transform 1 0 34684 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_370
timestamp 1667941163
transform 1 0 35144 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_374
timestamp 1667941163
transform 1 0 35512 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_380
timestamp 1667941163
transform 1 0 36064 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_402
timestamp 1667941163
transform 1 0 38088 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1667941163
transform 1 0 38456 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1667941163
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1667941163
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1667941163
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1667941163
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1667941163
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1667941163
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1667941163
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1667941163
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1667941163
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1667941163
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1667941163
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1667941163
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1667941163
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1667941163
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1667941163
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1667941163
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1667941163
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1667941163
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_169
timestamp 1667941163
transform 1 0 16652 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_179
timestamp 1667941163
transform 1 0 17572 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_194
timestamp 1667941163
transform 1 0 18952 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_208
timestamp 1667941163
transform 1 0 20240 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_215
timestamp 1667941163
transform 1 0 20884 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1667941163
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_225
timestamp 1667941163
transform 1 0 21804 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_229
timestamp 1667941163
transform 1 0 22172 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_236
timestamp 1667941163
transform 1 0 22816 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_245
timestamp 1667941163
transform 1 0 23644 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_258
timestamp 1667941163
transform 1 0 24840 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_266
timestamp 1667941163
transform 1 0 25576 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1667941163
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_47_281
timestamp 1667941163
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_286
timestamp 1667941163
transform 1 0 27416 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_300
timestamp 1667941163
transform 1 0 28704 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_312
timestamp 1667941163
transform 1 0 29808 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_321
timestamp 1667941163
transform 1 0 30636 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1667941163
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1667941163
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_337
timestamp 1667941163
transform 1 0 32108 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_355
timestamp 1667941163
transform 1 0 33764 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_362
timestamp 1667941163
transform 1 0 34408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_369
timestamp 1667941163
transform 1 0 35052 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_377
timestamp 1667941163
transform 1 0 35788 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_382
timestamp 1667941163
transform 1 0 36248 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_47_389
timestamp 1667941163
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_393
timestamp 1667941163
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_47_400
timestamp 1667941163
transform 1 0 37904 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_406
timestamp 1667941163
transform 1 0 38456 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1667941163
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1667941163
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1667941163
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1667941163
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1667941163
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1667941163
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1667941163
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1667941163
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1667941163
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1667941163
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1667941163
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1667941163
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1667941163
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1667941163
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1667941163
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1667941163
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1667941163
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1667941163
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1667941163
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1667941163
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1667941163
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_197
timestamp 1667941163
transform 1 0 19228 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_219
timestamp 1667941163
transform 1 0 21252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_231
timestamp 1667941163
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_240
timestamp 1667941163
transform 1 0 23184 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1667941163
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_253
timestamp 1667941163
transform 1 0 24380 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_259
timestamp 1667941163
transform 1 0 24932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_48_276
timestamp 1667941163
transform 1 0 26496 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_48_288
timestamp 1667941163
transform 1 0 27600 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_300
timestamp 1667941163
transform 1 0 28704 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1667941163
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_316
timestamp 1667941163
transform 1 0 30176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_325
timestamp 1667941163
transform 1 0 31004 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_345
timestamp 1667941163
transform 1 0 32844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_352
timestamp 1667941163
transform 1 0 33488 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_48_361
timestamp 1667941163
transform 1 0 34316 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_365
timestamp 1667941163
transform 1 0 34684 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_383
timestamp 1667941163
transform 1 0 36340 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1667941163
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1667941163
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1667941163
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1667941163
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1667941163
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1667941163
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1667941163
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1667941163
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1667941163
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1667941163
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1667941163
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1667941163
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1667941163
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1667941163
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1667941163
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1667941163
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1667941163
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1667941163
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1667941163
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_169
timestamp 1667941163
transform 1 0 16652 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_49_178
timestamp 1667941163
transform 1 0 17480 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_190
timestamp 1667941163
transform 1 0 18584 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_194
timestamp 1667941163
transform 1 0 18952 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_206
timestamp 1667941163
transform 1 0 20056 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1667941163
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1667941163
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_232
timestamp 1667941163
transform 1 0 22448 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_252
timestamp 1667941163
transform 1 0 24288 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_264
timestamp 1667941163
transform 1 0 25392 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_271
timestamp 1667941163
transform 1 0 26036 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1667941163
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_281
timestamp 1667941163
transform 1 0 26956 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_289
timestamp 1667941163
transform 1 0 27692 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_297
timestamp 1667941163
transform 1 0 28428 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_304
timestamp 1667941163
transform 1 0 29072 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_308
timestamp 1667941163
transform 1 0 29440 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_325
timestamp 1667941163
transform 1 0 31004 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_49_334
timestamp 1667941163
transform 1 0 31832 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_337
timestamp 1667941163
transform 1 0 32108 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_348
timestamp 1667941163
transform 1 0 33120 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_354
timestamp 1667941163
transform 1 0 33672 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_361
timestamp 1667941163
transform 1 0 34316 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_369
timestamp 1667941163
transform 1 0 35052 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_376
timestamp 1667941163
transform 1 0 35696 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_382
timestamp 1667941163
transform 1 0 36248 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_388
timestamp 1667941163
transform 1 0 36800 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_393
timestamp 1667941163
transform 1 0 37260 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_49_400
timestamp 1667941163
transform 1 0 37904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_406
timestamp 1667941163
transform 1 0 38456 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1667941163
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1667941163
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1667941163
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1667941163
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1667941163
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1667941163
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1667941163
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1667941163
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1667941163
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1667941163
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1667941163
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1667941163
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1667941163
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1667941163
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1667941163
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1667941163
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1667941163
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_165
timestamp 1667941163
transform 1 0 16284 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_169
timestamp 1667941163
transform 1 0 16652 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_180
timestamp 1667941163
transform 1 0 17664 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_188
timestamp 1667941163
transform 1 0 18400 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_194
timestamp 1667941163
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1667941163
transform 1 0 19228 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_50_207
timestamp 1667941163
transform 1 0 20148 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_215
timestamp 1667941163
transform 1 0 20884 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_220
timestamp 1667941163
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_233
timestamp 1667941163
transform 1 0 22540 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1667941163
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1667941163
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_253
timestamp 1667941163
transform 1 0 24380 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_261
timestamp 1667941163
transform 1 0 25116 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_265
timestamp 1667941163
transform 1 0 25484 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_272
timestamp 1667941163
transform 1 0 26128 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_50_286
timestamp 1667941163
transform 1 0 27416 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_294
timestamp 1667941163
transform 1 0 28152 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1667941163
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_309
timestamp 1667941163
transform 1 0 29532 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_318
timestamp 1667941163
transform 1 0 30360 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_330
timestamp 1667941163
transform 1 0 31464 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_50_338
timestamp 1667941163
transform 1 0 32200 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_350
timestamp 1667941163
transform 1 0 33304 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_354
timestamp 1667941163
transform 1 0 33672 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_362
timestamp 1667941163
transform 1 0 34408 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_365
timestamp 1667941163
transform 1 0 34684 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_50_372
timestamp 1667941163
transform 1 0 35328 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_378
timestamp 1667941163
transform 1 0 35880 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_385
timestamp 1667941163
transform 1 0 36524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_405
timestamp 1667941163
transform 1 0 38364 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1667941163
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1667941163
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1667941163
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1667941163
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1667941163
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1667941163
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1667941163
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1667941163
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1667941163
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1667941163
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1667941163
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1667941163
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1667941163
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1667941163
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1667941163
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1667941163
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1667941163
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1667941163
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_51_169
timestamp 1667941163
transform 1 0 16652 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_175
timestamp 1667941163
transform 1 0 17204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_186
timestamp 1667941163
transform 1 0 18216 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1667941163
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_219
timestamp 1667941163
transform 1 0 21252 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1667941163
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_225
timestamp 1667941163
transform 1 0 21804 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_51_237
timestamp 1667941163
transform 1 0 22908 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_243
timestamp 1667941163
transform 1 0 23460 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_260
timestamp 1667941163
transform 1 0 25024 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_271
timestamp 1667941163
transform 1 0 26036 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1667941163
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_281
timestamp 1667941163
transform 1 0 26956 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_299
timestamp 1667941163
transform 1 0 28612 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_311
timestamp 1667941163
transform 1 0 29716 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_323
timestamp 1667941163
transform 1 0 30820 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1667941163
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1667941163
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_349
timestamp 1667941163
transform 1 0 33212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_51_365
timestamp 1667941163
transform 1 0 34684 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_371
timestamp 1667941163
transform 1 0 35236 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_388
timestamp 1667941163
transform 1 0 36800 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_393
timestamp 1667941163
transform 1 0 37260 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_402
timestamp 1667941163
transform 1 0 38088 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_406
timestamp 1667941163
transform 1 0 38456 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_3
timestamp 1667941163
transform 1 0 1380 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_9
timestamp 1667941163
transform 1 0 1932 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_21
timestamp 1667941163
transform 1 0 3036 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1667941163
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1667941163
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1667941163
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1667941163
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1667941163
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1667941163
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1667941163
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1667941163
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1667941163
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1667941163
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1667941163
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1667941163
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1667941163
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1667941163
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1667941163
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_165
timestamp 1667941163
transform 1 0 16284 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_179
timestamp 1667941163
transform 1 0 17572 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1667941163
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1667941163
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_197
timestamp 1667941163
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_204
timestamp 1667941163
transform 1 0 19872 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_211
timestamp 1667941163
transform 1 0 20516 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_219
timestamp 1667941163
transform 1 0 21252 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_237
timestamp 1667941163
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_249
timestamp 1667941163
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_253
timestamp 1667941163
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_52_258
timestamp 1667941163
transform 1 0 24840 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_264
timestamp 1667941163
transform 1 0 25392 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_269
timestamp 1667941163
transform 1 0 25852 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_276
timestamp 1667941163
transform 1 0 26496 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_283
timestamp 1667941163
transform 1 0 27140 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_295
timestamp 1667941163
transform 1 0 28244 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_301
timestamp 1667941163
transform 1 0 28796 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_306
timestamp 1667941163
transform 1 0 29256 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_309
timestamp 1667941163
transform 1 0 29532 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_317
timestamp 1667941163
transform 1 0 30268 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_341
timestamp 1667941163
transform 1 0 32476 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1667941163
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_52_365
timestamp 1667941163
transform 1 0 34684 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_371
timestamp 1667941163
transform 1 0 35236 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_375
timestamp 1667941163
transform 1 0 35604 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_384
timestamp 1667941163
transform 1 0 36432 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_388
timestamp 1667941163
transform 1 0 36800 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_52_405
timestamp 1667941163
transform 1 0 38364 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1667941163
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1667941163
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1667941163
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1667941163
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1667941163
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1667941163
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1667941163
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1667941163
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1667941163
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1667941163
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1667941163
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1667941163
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1667941163
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1667941163
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1667941163
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1667941163
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1667941163
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1667941163
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1667941163
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1667941163
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_193
timestamp 1667941163
transform 1 0 18860 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_199
timestamp 1667941163
transform 1 0 19412 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_53_216
timestamp 1667941163
transform 1 0 20976 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_225
timestamp 1667941163
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_53_233
timestamp 1667941163
transform 1 0 22540 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_245
timestamp 1667941163
transform 1 0 23644 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_257
timestamp 1667941163
transform 1 0 24748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_269
timestamp 1667941163
transform 1 0 25852 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_277
timestamp 1667941163
transform 1 0 26588 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_53_281
timestamp 1667941163
transform 1 0 26956 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_289
timestamp 1667941163
transform 1 0 27692 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_306
timestamp 1667941163
transform 1 0 29256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_326
timestamp 1667941163
transform 1 0 31096 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_53_333
timestamp 1667941163
transform 1 0 31740 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_53_337
timestamp 1667941163
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_343
timestamp 1667941163
transform 1 0 32660 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_352
timestamp 1667941163
transform 1 0 33488 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_364
timestamp 1667941163
transform 1 0 34592 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_372
timestamp 1667941163
transform 1 0 35328 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_390
timestamp 1667941163
transform 1 0 36984 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_393
timestamp 1667941163
transform 1 0 37260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_400
timestamp 1667941163
transform 1 0 37904 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_406
timestamp 1667941163
transform 1 0 38456 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1667941163
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1667941163
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1667941163
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1667941163
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1667941163
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1667941163
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1667941163
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1667941163
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1667941163
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1667941163
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1667941163
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1667941163
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1667941163
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1667941163
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1667941163
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1667941163
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1667941163
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1667941163
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1667941163
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1667941163
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1667941163
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1667941163
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_209
timestamp 1667941163
transform 1 0 20332 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_54_217
timestamp 1667941163
transform 1 0 21068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_224
timestamp 1667941163
transform 1 0 21712 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_244
timestamp 1667941163
transform 1 0 23552 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_253
timestamp 1667941163
transform 1 0 24380 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_263
timestamp 1667941163
transform 1 0 25300 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_287
timestamp 1667941163
transform 1 0 27508 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_299
timestamp 1667941163
transform 1 0 28612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1667941163
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_309
timestamp 1667941163
transform 1 0 29532 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_54_315
timestamp 1667941163
transform 1 0 30084 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_337
timestamp 1667941163
transform 1 0 32108 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1667941163
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1667941163
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_365
timestamp 1667941163
transform 1 0 34684 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_383
timestamp 1667941163
transform 1 0 36340 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_390
timestamp 1667941163
transform 1 0 36984 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_394
timestamp 1667941163
transform 1 0 37352 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_398
timestamp 1667941163
transform 1 0 37720 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_54_405
timestamp 1667941163
transform 1 0 38364 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1667941163
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1667941163
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1667941163
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1667941163
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1667941163
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1667941163
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1667941163
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1667941163
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1667941163
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1667941163
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1667941163
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1667941163
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1667941163
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1667941163
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1667941163
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1667941163
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1667941163
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1667941163
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1667941163
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1667941163
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1667941163
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1667941163
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1667941163
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1667941163
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1667941163
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_237
timestamp 1667941163
transform 1 0 22908 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_252
timestamp 1667941163
transform 1 0 24288 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_263
timestamp 1667941163
transform 1 0 25300 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_271
timestamp 1667941163
transform 1 0 26036 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1667941163
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_281
timestamp 1667941163
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_289
timestamp 1667941163
transform 1 0 27692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_300
timestamp 1667941163
transform 1 0 28704 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_307
timestamp 1667941163
transform 1 0 29348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_315
timestamp 1667941163
transform 1 0 30084 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_325
timestamp 1667941163
transform 1 0 31004 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_333
timestamp 1667941163
transform 1 0 31740 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1667941163
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_349
timestamp 1667941163
transform 1 0 33212 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_358
timestamp 1667941163
transform 1 0 34040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_367
timestamp 1667941163
transform 1 0 34868 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_374
timestamp 1667941163
transform 1 0 35512 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_386
timestamp 1667941163
transform 1 0 36616 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_393
timestamp 1667941163
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_398
timestamp 1667941163
transform 1 0 37720 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_406
timestamp 1667941163
transform 1 0 38456 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1667941163
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1667941163
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1667941163
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1667941163
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1667941163
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1667941163
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1667941163
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1667941163
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1667941163
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1667941163
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1667941163
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1667941163
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1667941163
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1667941163
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1667941163
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1667941163
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1667941163
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1667941163
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1667941163
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1667941163
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1667941163
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1667941163
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1667941163
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1667941163
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_233
timestamp 1667941163
transform 1 0 22540 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_237
timestamp 1667941163
transform 1 0 22908 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_242
timestamp 1667941163
transform 1 0 23368 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_250
timestamp 1667941163
transform 1 0 24104 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_253
timestamp 1667941163
transform 1 0 24380 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_56_266
timestamp 1667941163
transform 1 0 25576 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_274
timestamp 1667941163
transform 1 0 26312 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_282
timestamp 1667941163
transform 1 0 27048 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_286
timestamp 1667941163
transform 1 0 27416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_291
timestamp 1667941163
transform 1 0 27876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_299
timestamp 1667941163
transform 1 0 28612 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_306
timestamp 1667941163
transform 1 0 29256 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_56_309
timestamp 1667941163
transform 1 0 29532 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_317
timestamp 1667941163
transform 1 0 30268 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_323
timestamp 1667941163
transform 1 0 30820 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_331
timestamp 1667941163
transform 1 0 31556 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_343
timestamp 1667941163
transform 1 0 32660 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_359
timestamp 1667941163
transform 1 0 34132 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1667941163
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_365
timestamp 1667941163
transform 1 0 34684 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_373
timestamp 1667941163
transform 1 0 35420 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_385
timestamp 1667941163
transform 1 0 36524 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_397
timestamp 1667941163
transform 1 0 37628 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_405
timestamp 1667941163
transform 1 0 38364 0 1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1667941163
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1667941163
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1667941163
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1667941163
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1667941163
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1667941163
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1667941163
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1667941163
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1667941163
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1667941163
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1667941163
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1667941163
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1667941163
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1667941163
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1667941163
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1667941163
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1667941163
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1667941163
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1667941163
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1667941163
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1667941163
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1667941163
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1667941163
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1667941163
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1667941163
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_237
timestamp 1667941163
transform 1 0 22908 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_57_252
timestamp 1667941163
transform 1 0 24288 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_261
timestamp 1667941163
transform 1 0 25116 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_269
timestamp 1667941163
transform 1 0 25852 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1667941163
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_281
timestamp 1667941163
transform 1 0 26956 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_290
timestamp 1667941163
transform 1 0 27784 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_301
timestamp 1667941163
transform 1 0 28796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_311
timestamp 1667941163
transform 1 0 29716 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_321
timestamp 1667941163
transform 1 0 30636 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1667941163
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1667941163
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_349
timestamp 1667941163
transform 1 0 33212 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_358
timestamp 1667941163
transform 1 0 34040 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_370
timestamp 1667941163
transform 1 0 35144 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1667941163
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1667941163
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1667941163
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1667941163
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1667941163
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1667941163
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1667941163
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1667941163
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1667941163
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1667941163
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1667941163
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1667941163
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1667941163
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1667941163
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1667941163
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1667941163
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1667941163
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1667941163
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1667941163
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1667941163
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1667941163
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1667941163
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1667941163
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1667941163
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1667941163
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1667941163
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1667941163
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1667941163
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1667941163
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1667941163
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1667941163
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_253
timestamp 1667941163
transform 1 0 24380 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_258
timestamp 1667941163
transform 1 0 24840 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_270
timestamp 1667941163
transform 1 0 25944 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_58_280
timestamp 1667941163
transform 1 0 26864 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_292
timestamp 1667941163
transform 1 0 27968 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_299
timestamp 1667941163
transform 1 0 28612 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1667941163
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_58_309
timestamp 1667941163
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1667941163
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_328
timestamp 1667941163
transform 1 0 31280 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_340
timestamp 1667941163
transform 1 0 32384 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_352
timestamp 1667941163
transform 1 0 33488 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1667941163
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1667941163
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1667941163
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1667941163
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1667941163
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1667941163
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1667941163
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1667941163
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1667941163
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1667941163
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1667941163
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1667941163
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1667941163
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1667941163
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1667941163
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1667941163
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1667941163
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1667941163
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1667941163
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1667941163
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1667941163
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1667941163
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1667941163
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1667941163
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1667941163
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1667941163
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1667941163
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1667941163
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1667941163
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1667941163
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1667941163
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1667941163
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1667941163
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1667941163
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1667941163
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1667941163
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1667941163
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1667941163
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1667941163
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1667941163
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1667941163
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1667941163
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1667941163
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1667941163
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1667941163
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1667941163
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1667941163
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1667941163
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1667941163
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1667941163
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1667941163
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1667941163
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1667941163
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1667941163
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1667941163
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1667941163
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1667941163
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1667941163
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1667941163
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1667941163
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1667941163
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1667941163
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1667941163
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1667941163
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1667941163
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1667941163
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1667941163
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1667941163
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1667941163
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1667941163
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1667941163
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1667941163
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1667941163
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1667941163
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1667941163
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1667941163
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1667941163
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1667941163
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1667941163
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1667941163
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1667941163
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1667941163
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1667941163
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1667941163
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1667941163
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1667941163
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1667941163
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1667941163
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1667941163
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1667941163
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1667941163
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1667941163
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1667941163
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1667941163
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1667941163
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1667941163
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1667941163
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1667941163
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1667941163
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_81
timestamp 1667941163
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_93
timestamp 1667941163
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_105
timestamp 1667941163
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1667941163
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1667941163
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1667941163
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1667941163
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1667941163
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1667941163
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1667941163
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1667941163
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1667941163
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1667941163
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1667941163
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1667941163
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1667941163
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1667941163
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1667941163
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1667941163
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1667941163
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1667941163
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1667941163
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1667941163
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1667941163
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1667941163
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1667941163
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1667941163
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1667941163
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1667941163
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1667941163
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1667941163
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1667941163
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1667941163
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1667941163
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1667941163
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1667941163
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1667941163
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1667941163
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1667941163
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1667941163
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1667941163
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1667941163
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1667941163
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1667941163
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1667941163
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1667941163
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1667941163
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1667941163
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1667941163
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1667941163
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1667941163
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1667941163
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1667941163
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1667941163
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1667941163
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1667941163
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1667941163
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1667941163
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1667941163
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1667941163
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1667941163
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1667941163
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1667941163
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1667941163
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1667941163
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1667941163
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1667941163
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1667941163
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1667941163
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1667941163
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1667941163
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1667941163
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1667941163
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1667941163
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1667941163
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1667941163
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1667941163
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1667941163
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1667941163
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1667941163
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1667941163
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1667941163
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1667941163
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1667941163
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1667941163
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1667941163
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1667941163
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1667941163
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1667941163
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1667941163
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1667941163
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1667941163
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1667941163
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1667941163
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1667941163
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1667941163
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1667941163
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1667941163
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1667941163
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1667941163
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1667941163
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1667941163
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1667941163
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1667941163
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1667941163
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1667941163
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1667941163
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1667941163
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1667941163
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1667941163
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1667941163
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1667941163
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1667941163
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1667941163
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1667941163
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_337
timestamp 1667941163
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_342
timestamp 1667941163
transform 1 0 32568 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_354
timestamp 1667941163
transform 1 0 33672 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_366
timestamp 1667941163
transform 1 0 34776 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_378
timestamp 1667941163
transform 1 0 35880 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_390
timestamp 1667941163
transform 1 0 36984 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1667941163
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1667941163
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_3
timestamp 1667941163
transform 1 0 1380 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_8
timestamp 1667941163
transform 1 0 1840 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_20
timestamp 1667941163
transform 1 0 2944 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1667941163
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1667941163
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1667941163
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1667941163
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1667941163
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1667941163
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1667941163
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_97
timestamp 1667941163
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_107
timestamp 1667941163
transform 1 0 10948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_111
timestamp 1667941163
transform 1 0 11316 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1667941163
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1667941163
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1667941163
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1667941163
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1667941163
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_165
timestamp 1667941163
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1667941163
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1667941163
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1667941163
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_197
timestamp 1667941163
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1667941163
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1667941163
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1667941163
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1667941163
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1667941163
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1667941163
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1667941163
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1667941163
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1667941163
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1667941163
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1667941163
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1667941163
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_64_309
timestamp 1667941163
transform 1 0 29532 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_314
timestamp 1667941163
transform 1 0 29992 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_326
timestamp 1667941163
transform 1 0 31096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1667941163
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1667941163
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1667941163
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1667941163
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1667941163
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1667941163
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1667941163
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_393
timestamp 1667941163
transform 1 0 37260 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1667941163
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1667941163
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1667941163
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1667941163
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1667941163
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1667941163
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1667941163
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1667941163
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1667941163
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1667941163
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1667941163
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1667941163
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1667941163
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1667941163
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1667941163
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1667941163
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1667941163
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1667941163
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1667941163
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1667941163
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1667941163
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1667941163
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1667941163
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1667941163
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1667941163
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1667941163
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1667941163
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1667941163
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1667941163
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1667941163
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1667941163
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1667941163
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1667941163
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1667941163
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1667941163
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1667941163
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1667941163
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1667941163
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1667941163
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1667941163
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1667941163
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1667941163
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1667941163
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1667941163
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1667941163
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1667941163
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1667941163
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1667941163
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1667941163
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1667941163
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1667941163
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1667941163
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1667941163
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1667941163
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1667941163
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1667941163
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1667941163
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1667941163
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1667941163
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1667941163
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1667941163
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1667941163
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1667941163
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1667941163
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1667941163
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1667941163
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1667941163
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1667941163
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1667941163
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1667941163
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1667941163
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1667941163
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1667941163
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1667941163
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1667941163
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1667941163
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1667941163
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1667941163
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1667941163
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1667941163
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1667941163
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1667941163
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1667941163
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1667941163
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1667941163
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1667941163
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1667941163
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1667941163
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1667941163
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1667941163
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1667941163
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1667941163
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1667941163
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1667941163
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1667941163
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1667941163
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1667941163
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1667941163
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1667941163
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1667941163
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1667941163
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1667941163
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1667941163
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1667941163
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1667941163
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1667941163
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1667941163
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1667941163
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1667941163
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1667941163
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1667941163
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1667941163
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1667941163
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1667941163
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1667941163
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1667941163
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1667941163
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1667941163
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1667941163
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1667941163
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1667941163
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1667941163
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1667941163
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1667941163
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1667941163
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1667941163
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1667941163
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1667941163
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1667941163
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1667941163
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1667941163
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1667941163
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1667941163
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1667941163
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1667941163
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1667941163
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1667941163
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1667941163
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1667941163
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1667941163
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1667941163
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1667941163
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1667941163
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1667941163
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1667941163
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1667941163
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1667941163
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1667941163
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1667941163
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1667941163
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1667941163
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1667941163
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1667941163
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1667941163
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1667941163
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1667941163
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1667941163
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1667941163
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1667941163
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1667941163
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1667941163
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1667941163
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1667941163
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1667941163
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1667941163
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1667941163
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1667941163
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1667941163
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1667941163
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1667941163
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1667941163
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1667941163
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1667941163
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1667941163
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1667941163
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1667941163
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1667941163
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1667941163
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1667941163
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1667941163
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1667941163
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1667941163
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1667941163
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1667941163
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1667941163
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1667941163
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1667941163
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1667941163
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1667941163
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1667941163
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1667941163
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1667941163
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1667941163
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1667941163
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1667941163
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1667941163
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1667941163
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1667941163
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1667941163
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1667941163
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1667941163
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1667941163
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1667941163
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1667941163
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1667941163
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1667941163
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1667941163
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1667941163
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1667941163
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1667941163
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1667941163
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1667941163
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1667941163
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1667941163
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1667941163
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1667941163
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1667941163
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1667941163
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1667941163
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1667941163
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1667941163
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1667941163
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1667941163
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1667941163
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1667941163
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1667941163
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1667941163
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1667941163
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1667941163
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1667941163
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1667941163
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1667941163
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1667941163
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1667941163
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1667941163
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1667941163
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1667941163
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1667941163
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1667941163
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1667941163
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1667941163
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1667941163
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1667941163
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1667941163
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1667941163
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1667941163
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1667941163
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1667941163
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1667941163
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1667941163
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1667941163
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1667941163
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1667941163
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1667941163
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1667941163
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1667941163
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1667941163
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1667941163
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1667941163
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1667941163
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1667941163
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1667941163
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1667941163
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1667941163
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1667941163
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1667941163
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1667941163
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1667941163
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1667941163
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1667941163
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1667941163
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1667941163
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1667941163
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1667941163
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1667941163
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1667941163
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1667941163
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1667941163
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1667941163
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1667941163
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1667941163
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1667941163
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1667941163
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1667941163
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1667941163
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1667941163
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1667941163
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1667941163
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1667941163
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1667941163
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1667941163
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1667941163
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1667941163
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1667941163
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1667941163
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1667941163
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1667941163
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1667941163
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1667941163
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1667941163
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1667941163
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1667941163
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1667941163
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1667941163
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1667941163
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1667941163
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1667941163
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1667941163
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1667941163
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1667941163
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1667941163
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1667941163
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1667941163
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1667941163
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1667941163
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1667941163
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1667941163
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1667941163
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1667941163
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1667941163
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1667941163
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1667941163
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1667941163
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1667941163
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1667941163
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1667941163
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1667941163
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1667941163
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1667941163
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1667941163
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1667941163
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1667941163
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1667941163
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1667941163
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1667941163
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1667941163
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1667941163
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1667941163
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1667941163
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1667941163
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1667941163
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1667941163
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1667941163
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1667941163
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1667941163
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1667941163
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1667941163
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1667941163
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1667941163
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1667941163
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1667941163
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1667941163
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1667941163
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1667941163
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1667941163
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1667941163
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1667941163
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1667941163
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1667941163
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1667941163
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1667941163
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1667941163
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1667941163
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1667941163
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1667941163
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1667941163
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1667941163
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1667941163
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1667941163
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1667941163
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1667941163
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1667941163
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1667941163
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1667941163
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1667941163
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1667941163
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1667941163
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1667941163
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1667941163
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1667941163
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1667941163
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1667941163
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1667941163
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1667941163
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1667941163
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1667941163
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1667941163
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1667941163
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1667941163
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1667941163
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1667941163
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1667941163
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1667941163
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1667941163
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1667941163
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1667941163
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1667941163
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1667941163
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1667941163
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1667941163
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1667941163
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1667941163
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1667941163
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1667941163
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1667941163
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1667941163
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1667941163
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1667941163
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1667941163
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1667941163
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1667941163
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1667941163
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1667941163
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1667941163
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1667941163
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1667941163
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1667941163
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1667941163
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1667941163
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1667941163
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1667941163
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1667941163
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1667941163
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1667941163
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1667941163
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1667941163
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1667941163
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1667941163
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1667941163
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1667941163
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1667941163
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1667941163
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1667941163
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1667941163
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1667941163
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1667941163
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1667941163
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1667941163
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1667941163
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1667941163
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1667941163
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1667941163
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1667941163
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1667941163
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1667941163
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1667941163
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1667941163
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1667941163
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1667941163
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1667941163
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1667941163
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1667941163
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1667941163
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1667941163
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1667941163
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1667941163
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1667941163
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1667941163
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1667941163
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1667941163
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1667941163
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1667941163
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1667941163
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1667941163
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1667941163
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1667941163
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1667941163
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1667941163
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1667941163
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1667941163
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1667941163
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1667941163
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1667941163
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1667941163
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1667941163
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1667941163
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1667941163
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1667941163
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1667941163
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1667941163
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1667941163
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1667941163
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1667941163
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1667941163
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1667941163
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1667941163
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1667941163
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1667941163
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1667941163
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1667941163
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1667941163
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1667941163
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1667941163
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1667941163
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1667941163
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1667941163
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1667941163
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1667941163
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1667941163
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1667941163
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1667941163
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1667941163
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1667941163
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1667941163
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1667941163
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1667941163
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1667941163
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1667941163
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1667941163
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1667941163
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1667941163
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1667941163
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1667941163
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1667941163
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1667941163
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1667941163
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1667941163
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1667941163
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1667941163
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1667941163
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1667941163
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1667941163
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1667941163
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1667941163
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1667941163
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1667941163
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1667941163
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1667941163
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1667941163
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1667941163
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1667941163
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1667941163
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1667941163
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1667941163
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1667941163
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1667941163
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1667941163
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1667941163
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1667941163
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1667941163
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1667941163
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1667941163
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1667941163
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1667941163
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1667941163
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1667941163
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1667941163
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1667941163
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1667941163
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1667941163
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1667941163
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1667941163
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1667941163
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1667941163
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1667941163
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1667941163
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1667941163
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1667941163
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1667941163
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1667941163
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1667941163
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1667941163
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1667941163
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1667941163
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1667941163
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1667941163
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1667941163
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1667941163
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1667941163
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1667941163
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1667941163
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1667941163
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1667941163
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1667941163
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1667941163
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1667941163
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1667941163
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1667941163
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1667941163
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1667941163
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1667941163
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1667941163
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1667941163
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1667941163
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1667941163
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1667941163
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1667941163
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1667941163
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1667941163
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1667941163
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1667941163
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1667941163
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1667941163
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1667941163
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1667941163
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1667941163
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1667941163
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1667941163
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1667941163
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_2  _426_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29532 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _427_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _428_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31004 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _429_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29900 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _430_
timestamp 1667941163
transform 1 0 32292 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1667941163
transform 1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _432_
timestamp 1667941163
transform 1 0 27968 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _433_
timestamp 1667941163
transform 1 0 27324 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _434_
timestamp 1667941163
transform 1 0 27140 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _435_
timestamp 1667941163
transform 1 0 26404 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _436_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27784 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _437_
timestamp 1667941163
transform 1 0 27140 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _438_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27968 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _439_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27968 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _440_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 26496 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _441_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27048 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _442_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 27508 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _443_
timestamp 1667941163
transform 1 0 28152 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _444_
timestamp 1667941163
transform 1 0 29716 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _445_
timestamp 1667941163
transform 1 0 29900 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _446_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30544 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _447_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32292 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1667941163
transform 1 0 20424 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _449_
timestamp 1667941163
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _450_
timestamp 1667941163
transform 1 0 22080 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _451_
timestamp 1667941163
transform 1 0 23552 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1667941163
transform 1 0 25760 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _453_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22724 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _454_
timestamp 1667941163
transform 1 0 26404 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _455_
timestamp 1667941163
transform 1 0 28060 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _456_
timestamp 1667941163
transform 1 0 28980 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _457_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 25484 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _458_
timestamp 1667941163
transform 1 0 24932 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _459_
timestamp 1667941163
transform 1 0 24656 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _460_
timestamp 1667941163
transform 1 0 23184 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _461_
timestamp 1667941163
transform 1 0 21988 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _462_
timestamp 1667941163
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _463_
timestamp 1667941163
transform 1 0 20240 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  _464_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19596 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _465_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 19596 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _466_
timestamp 1667941163
transform 1 0 20240 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _467_
timestamp 1667941163
transform 1 0 21068 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _468_
timestamp 1667941163
transform 1 0 21252 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _469_
timestamp 1667941163
transform 1 0 21252 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _470_
timestamp 1667941163
transform 1 0 22816 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _471_
timestamp 1667941163
transform 1 0 21988 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _472_
timestamp 1667941163
transform 1 0 20976 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _473_
timestamp 1667941163
transform 1 0 21252 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _474_
timestamp 1667941163
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _475_
timestamp 1667941163
transform 1 0 21344 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _476_
timestamp 1667941163
transform 1 0 21988 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _477_
timestamp 1667941163
transform 1 0 21620 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _478_
timestamp 1667941163
transform 1 0 21620 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _479_
timestamp 1667941163
transform 1 0 21988 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _480_
timestamp 1667941163
transform 1 0 21620 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _481_
timestamp 1667941163
transform 1 0 21712 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_2  _482_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 21988 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _483_
timestamp 1667941163
transform 1 0 33028 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _484_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 37444 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _485_
timestamp 1667941163
transform 1 0 33764 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _486_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _487_
timestamp 1667941163
transform 1 0 35972 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _488_
timestamp 1667941163
transform 1 0 34868 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _489_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33948 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _490_
timestamp 1667941163
transform 1 0 34132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _491_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33948 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _492_
timestamp 1667941163
transform 1 0 32384 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _493_
timestamp 1667941163
transform 1 0 21252 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _494_
timestamp 1667941163
transform 1 0 31464 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _495_
timestamp 1667941163
transform 1 0 31740 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _496_
timestamp 1667941163
transform 1 0 31556 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _497_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31464 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _498_
timestamp 1667941163
transform 1 0 32660 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _499_
timestamp 1667941163
transform 1 0 33212 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _500_
timestamp 1667941163
transform 1 0 33856 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _501_
timestamp 1667941163
transform 1 0 34776 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _502_
timestamp 1667941163
transform 1 0 35236 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _503_
timestamp 1667941163
transform 1 0 35328 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _504_
timestamp 1667941163
transform 1 0 35972 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _505_
timestamp 1667941163
transform 1 0 36708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _506_
timestamp 1667941163
transform 1 0 37444 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _507_
timestamp 1667941163
transform 1 0 37444 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _508_
timestamp 1667941163
transform 1 0 37444 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _509_
timestamp 1667941163
transform 1 0 37444 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _510_
timestamp 1667941163
transform 1 0 33488 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _511_
timestamp 1667941163
transform 1 0 34868 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _512_
timestamp 1667941163
transform 1 0 37444 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _513_
timestamp 1667941163
transform 1 0 36064 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _514_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 35604 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _515_
timestamp 1667941163
transform 1 0 36432 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _516_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 36156 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _517_
timestamp 1667941163
transform 1 0 34868 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _518_
timestamp 1667941163
transform 1 0 36340 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _519_
timestamp 1667941163
transform 1 0 35972 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _520_
timestamp 1667941163
transform 1 0 37444 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _521_
timestamp 1667941163
transform 1 0 36616 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _522_
timestamp 1667941163
transform 1 0 37444 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _523_
timestamp 1667941163
transform 1 0 36064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _524_
timestamp 1667941163
transform 1 0 34776 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _525_
timestamp 1667941163
transform 1 0 34868 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _526_
timestamp 1667941163
transform 1 0 37444 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _527_
timestamp 1667941163
transform 1 0 36708 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _528_
timestamp 1667941163
transform 1 0 33396 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _529_
timestamp 1667941163
transform 1 0 37444 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _530_
timestamp 1667941163
transform 1 0 37352 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _531_
timestamp 1667941163
transform 1 0 37444 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _532_
timestamp 1667941163
transform 1 0 36616 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _533_
timestamp 1667941163
transform 1 0 34868 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _534_
timestamp 1667941163
transform 1 0 34500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _535_
timestamp 1667941163
transform 1 0 36340 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _536_
timestamp 1667941163
transform 1 0 37444 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _537_
timestamp 1667941163
transform 1 0 36432 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _538_
timestamp 1667941163
transform 1 0 36340 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _539_
timestamp 1667941163
transform 1 0 35236 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _540_
timestamp 1667941163
transform 1 0 34408 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _541_
timestamp 1667941163
transform 1 0 35788 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _542_
timestamp 1667941163
transform 1 0 35236 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _543_
timestamp 1667941163
transform 1 0 35604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _544_
timestamp 1667941163
transform 1 0 35788 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _545_
timestamp 1667941163
transform 1 0 36524 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _546_
timestamp 1667941163
transform 1 0 37444 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _547_
timestamp 1667941163
transform 1 0 37352 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _548_
timestamp 1667941163
transform 1 0 37444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _549_
timestamp 1667941163
transform 1 0 37444 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _550_
timestamp 1667941163
transform 1 0 38088 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _551_
timestamp 1667941163
transform 1 0 36064 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _552_
timestamp 1667941163
transform 1 0 37444 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _553_
timestamp 1667941163
transform 1 0 35420 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _554_
timestamp 1667941163
transform 1 0 35236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _555_
timestamp 1667941163
transform 1 0 33396 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _556_
timestamp 1667941163
transform 1 0 33488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _557_
timestamp 1667941163
transform 1 0 34960 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _558_
timestamp 1667941163
transform 1 0 33856 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _559_
timestamp 1667941163
transform 1 0 32568 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _560_
timestamp 1667941163
transform 1 0 35972 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _561_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32752 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _562_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32568 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _563_
timestamp 1667941163
transform 1 0 24380 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _564_
timestamp 1667941163
transform 1 0 28980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _565_
timestamp 1667941163
transform 1 0 33120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _566_
timestamp 1667941163
transform 1 0 30544 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _567_
timestamp 1667941163
transform 1 0 31372 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _568_
timestamp 1667941163
transform 1 0 31924 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _569_
timestamp 1667941163
transform 1 0 31464 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _570_
timestamp 1667941163
transform 1 0 33856 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _571_
timestamp 1667941163
transform 1 0 34868 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _572_
timestamp 1667941163
transform 1 0 33948 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _573_
timestamp 1667941163
transform 1 0 34224 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 1667941163
transform 1 0 34408 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _575_
timestamp 1667941163
transform 1 0 35972 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _576_
timestamp 1667941163
transform 1 0 35144 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _577_
timestamp 1667941163
transform 1 0 36616 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _578_
timestamp 1667941163
transform 1 0 29992 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _579_
timestamp 1667941163
transform 1 0 28244 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _580_
timestamp 1667941163
transform 1 0 28244 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _581_
timestamp 1667941163
transform 1 0 28152 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _582_
timestamp 1667941163
transform 1 0 28244 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _583_
timestamp 1667941163
transform 1 0 31096 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _584_
timestamp 1667941163
transform 1 0 28980 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _585_
timestamp 1667941163
transform 1 0 27692 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _586_
timestamp 1667941163
transform 1 0 27968 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _587_
timestamp 1667941163
transform 1 0 22172 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _588_
timestamp 1667941163
transform 1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _589_
timestamp 1667941163
transform 1 0 25852 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _590_
timestamp 1667941163
transform 1 0 25668 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _591_
timestamp 1667941163
transform 1 0 27140 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _592_
timestamp 1667941163
transform 1 0 26404 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _593_
timestamp 1667941163
transform 1 0 28980 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _594_
timestamp 1667941163
transform 1 0 28336 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _595_
timestamp 1667941163
transform 1 0 29716 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _596_
timestamp 1667941163
transform 1 0 29256 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _597_
timestamp 1667941163
transform 1 0 30912 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _598_
timestamp 1667941163
transform 1 0 28704 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _599_
timestamp 1667941163
transform 1 0 28336 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _600_
timestamp 1667941163
transform 1 0 27416 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _601_
timestamp 1667941163
transform 1 0 29716 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _602_
timestamp 1667941163
transform 1 0 26588 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _603_
timestamp 1667941163
transform 1 0 27140 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _604_
timestamp 1667941163
transform 1 0 33212 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _605_
timestamp 1667941163
transform 1 0 34040 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _606_
timestamp 1667941163
transform 1 0 32292 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _607_
timestamp 1667941163
transform 1 0 33212 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _608_
timestamp 1667941163
transform 1 0 32292 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _609_
timestamp 1667941163
transform 1 0 32292 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _610_
timestamp 1667941163
transform 1 0 32292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _611_
timestamp 1667941163
transform 1 0 32108 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _612_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23828 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _613_
timestamp 1667941163
transform 1 0 24656 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _614_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23000 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _615_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 22080 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _616_
timestamp 1667941163
transform 1 0 23736 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _617_
timestamp 1667941163
transform 1 0 22540 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _618_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _619_
timestamp 1667941163
transform 1 0 22908 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _620_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _621_
timestamp 1667941163
transform 1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _622_
timestamp 1667941163
transform 1 0 22540 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _623_
timestamp 1667941163
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _624_
timestamp 1667941163
transform 1 0 22908 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _625_
timestamp 1667941163
transform 1 0 23184 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _626_
timestamp 1667941163
transform 1 0 23552 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _627_
timestamp 1667941163
transform 1 0 22264 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _628_
timestamp 1667941163
transform 1 0 22724 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _629_
timestamp 1667941163
transform 1 0 23552 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _630_
timestamp 1667941163
transform 1 0 22172 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _631_
timestamp 1667941163
transform 1 0 22908 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _632_
timestamp 1667941163
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _633_
timestamp 1667941163
transform 1 0 29716 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _634_
timestamp 1667941163
transform 1 0 29992 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _635_
timestamp 1667941163
transform 1 0 31372 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _636_
timestamp 1667941163
transform 1 0 33396 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _637_
timestamp 1667941163
transform 1 0 30912 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _638_
timestamp 1667941163
transform 1 0 29532 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _639_
timestamp 1667941163
transform 1 0 31096 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _640_
timestamp 1667941163
transform 1 0 30728 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _641_
timestamp 1667941163
transform 1 0 30360 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _642_
timestamp 1667941163
transform 1 0 30544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _643_
timestamp 1667941163
transform 1 0 31372 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _644_
timestamp 1667941163
transform 1 0 30728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _645_
timestamp 1667941163
transform 1 0 33396 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _646_
timestamp 1667941163
transform 1 0 34040 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _647_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 34868 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _648_
timestamp 1667941163
transform 1 0 33488 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _649_
timestamp 1667941163
transform 1 0 34408 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _650_
timestamp 1667941163
transform 1 0 35236 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _651_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 33396 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _652_
timestamp 1667941163
transform 1 0 29716 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _653_
timestamp 1667941163
transform 1 0 28888 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _654_
timestamp 1667941163
transform 1 0 29716 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _655_
timestamp 1667941163
transform 1 0 33396 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _656_
timestamp 1667941163
transform 1 0 30360 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _657_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 31004 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _658_
timestamp 1667941163
transform 1 0 30268 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _659_
timestamp 1667941163
transform 1 0 31004 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _660_
timestamp 1667941163
transform 1 0 31188 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _661_
timestamp 1667941163
transform 1 0 30176 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _662_
timestamp 1667941163
transform 1 0 30268 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _663_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 30084 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _664_
timestamp 1667941163
transform 1 0 28796 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _665_
timestamp 1667941163
transform 1 0 29164 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _666_
timestamp 1667941163
transform 1 0 28336 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _667_
timestamp 1667941163
transform 1 0 28980 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _668_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28152 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _669_
timestamp 1667941163
transform 1 0 29072 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _670_
timestamp 1667941163
transform 1 0 27968 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _671_
timestamp 1667941163
transform 1 0 25944 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _672_
timestamp 1667941163
transform 1 0 27600 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21boi_1  _673_
timestamp 1667941163
transform 1 0 26496 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _674_
timestamp 1667941163
transform 1 0 26496 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _675_
timestamp 1667941163
transform 1 0 27876 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _676_
timestamp 1667941163
transform 1 0 27508 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _677_
timestamp 1667941163
transform 1 0 27140 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _678_
timestamp 1667941163
transform 1 0 23644 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _679_
timestamp 1667941163
transform 1 0 24656 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _680_
timestamp 1667941163
transform 1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _681_
timestamp 1667941163
transform 1 0 23000 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _682_
timestamp 1667941163
transform 1 0 24564 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _683_
timestamp 1667941163
transform 1 0 24656 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _684_
timestamp 1667941163
transform 1 0 23736 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _685_
timestamp 1667941163
transform 1 0 23644 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _686_
timestamp 1667941163
transform 1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _687_
timestamp 1667941163
transform 1 0 24564 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _688_
timestamp 1667941163
transform 1 0 26220 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _689_
timestamp 1667941163
transform 1 0 26404 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _690_
timestamp 1667941163
transform 1 0 25576 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _691_
timestamp 1667941163
transform 1 0 25668 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _692_
timestamp 1667941163
transform 1 0 24932 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _693_
timestamp 1667941163
transform 1 0 25392 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _694_
timestamp 1667941163
transform 1 0 26864 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _695_
timestamp 1667941163
transform 1 0 26680 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _696_
timestamp 1667941163
transform 1 0 25484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _697_
timestamp 1667941163
transform 1 0 29716 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _698_
timestamp 1667941163
transform 1 0 28796 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _699_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 28980 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _700_
timestamp 1667941163
transform 1 0 28428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _701_
timestamp 1667941163
transform 1 0 33764 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _702_
timestamp 1667941163
transform 1 0 34868 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _703_
timestamp 1667941163
transform 1 0 33028 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _704_
timestamp 1667941163
transform 1 0 32384 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _705_
timestamp 1667941163
transform 1 0 33856 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _706_
timestamp 1667941163
transform 1 0 33672 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _707_
timestamp 1667941163
transform 1 0 32752 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _708_
timestamp 1667941163
transform 1 0 33028 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _709_
timestamp 1667941163
transform 1 0 32660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _710_
timestamp 1667941163
transform 1 0 20976 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _711_
timestamp 1667941163
transform 1 0 27140 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _712_
timestamp 1667941163
transform 1 0 27140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _713_
timestamp 1667941163
transform 1 0 32660 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _714_
timestamp 1667941163
transform 1 0 28060 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _715_
timestamp 1667941163
transform 1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _716_
timestamp 1667941163
transform 1 0 27416 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _717_
timestamp 1667941163
transform 1 0 27416 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _718_
timestamp 1667941163
transform 1 0 26680 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _719_
timestamp 1667941163
transform 1 0 28428 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _720_
timestamp 1667941163
transform 1 0 27140 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _721_
timestamp 1667941163
transform 1 0 27692 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _722_
timestamp 1667941163
transform 1 0 27232 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _723_
timestamp 1667941163
transform 1 0 27232 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _724_
timestamp 1667941163
transform 1 0 28152 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _725_
timestamp 1667941163
transform 1 0 27416 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _726_
timestamp 1667941163
transform 1 0 28428 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _727_
timestamp 1667941163
transform 1 0 28520 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _728_
timestamp 1667941163
transform 1 0 25208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _729_
timestamp 1667941163
transform 1 0 26680 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _730_
timestamp 1667941163
transform 1 0 25576 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _731_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 24656 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _732_
timestamp 1667941163
transform 1 0 25116 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _733_
timestamp 1667941163
transform 1 0 26220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _734_
timestamp 1667941163
transform 1 0 25944 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _735_
timestamp 1667941163
transform 1 0 23460 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _736_
timestamp 1667941163
transform 1 0 23736 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _737_
timestamp 1667941163
transform 1 0 24564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _738_
timestamp 1667941163
transform 1 0 23736 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _739_
timestamp 1667941163
transform 1 0 23368 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _740_
timestamp 1667941163
transform 1 0 21988 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _741_
timestamp 1667941163
transform 1 0 23460 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _742_
timestamp 1667941163
transform 1 0 22264 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _743_
timestamp 1667941163
transform 1 0 22356 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _744_
timestamp 1667941163
transform 1 0 22172 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _745_
timestamp 1667941163
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _746_
timestamp 1667941163
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _747_
timestamp 1667941163
transform 1 0 20332 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _748_
timestamp 1667941163
transform 1 0 22908 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _749_
timestamp 1667941163
transform 1 0 23000 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _750_
timestamp 1667941163
transform 1 0 20332 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _751_
timestamp 1667941163
transform 1 0 21160 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _752_
timestamp 1667941163
transform 1 0 21252 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _753_
timestamp 1667941163
transform 1 0 20056 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _754_
timestamp 1667941163
transform 1 0 18676 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _755_
timestamp 1667941163
transform 1 0 19596 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _756_
timestamp 1667941163
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _757_
timestamp 1667941163
transform 1 0 19688 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _758_
timestamp 1667941163
transform 1 0 31372 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _759_
timestamp 1667941163
transform 1 0 30084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _760_
timestamp 1667941163
transform 1 0 26496 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _761_
timestamp 1667941163
transform 1 0 26128 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _762_
timestamp 1667941163
transform 1 0 24932 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _763_
timestamp 1667941163
transform 1 0 26864 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_2  _764_
timestamp 1667941163
transform 1 0 25760 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _765_
timestamp 1667941163
transform 1 0 19412 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _766_
timestamp 1667941163
transform 1 0 20976 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _767_
timestamp 1667941163
transform 1 0 20056 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _768_
timestamp 1667941163
transform 1 0 25760 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _769_
timestamp 1667941163
transform 1 0 18400 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _770_
timestamp 1667941163
transform 1 0 17756 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _771_
timestamp 1667941163
transform 1 0 17664 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _772_
timestamp 1667941163
transform 1 0 18400 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _773_
timestamp 1667941163
transform 1 0 18584 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _774_
timestamp 1667941163
transform 1 0 18492 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__a21boi_1  _775_
timestamp 1667941163
transform 1 0 17572 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _776_
timestamp 1667941163
transform 1 0 17756 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _777_
timestamp 1667941163
transform 1 0 17756 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _778_
timestamp 1667941163
transform 1 0 16100 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _779_
timestamp 1667941163
transform 1 0 18676 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _780_
timestamp 1667941163
transform 1 0 17664 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _781_
timestamp 1667941163
transform 1 0 19228 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _782_
timestamp 1667941163
transform 1 0 19504 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _783_
timestamp 1667941163
transform 1 0 17388 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _784_
timestamp 1667941163
transform 1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _785_
timestamp 1667941163
transform 1 0 18216 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21bai_1  _786_
timestamp 1667941163
transform 1 0 18584 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _787_
timestamp 1667941163
transform 1 0 19412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _788_
timestamp 1667941163
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _789_
timestamp 1667941163
transform 1 0 17204 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _790_
timestamp 1667941163
transform 1 0 16284 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _791_
timestamp 1667941163
transform 1 0 17756 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _792_
timestamp 1667941163
transform 1 0 17848 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _793_
timestamp 1667941163
transform 1 0 18492 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _794_
timestamp 1667941163
transform 1 0 18584 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _795_
timestamp 1667941163
transform 1 0 16928 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _796_
timestamp 1667941163
transform 1 0 18308 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _797_
timestamp 1667941163
transform 1 0 18308 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _798_
timestamp 1667941163
transform 1 0 20608 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _799_
timestamp 1667941163
transform 1 0 19688 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _800_
timestamp 1667941163
transform 1 0 16928 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _801_
timestamp 1667941163
transform 1 0 16376 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _802_
timestamp 1667941163
transform 1 0 17020 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _803_
timestamp 1667941163
transform 1 0 17020 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _804_
timestamp 1667941163
transform 1 0 17296 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _805_
timestamp 1667941163
transform 1 0 17020 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _806_
timestamp 1667941163
transform 1 0 18676 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _807_
timestamp 1667941163
transform 1 0 19412 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _808_
timestamp 1667941163
transform 1 0 16928 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _809_
timestamp 1667941163
transform 1 0 17572 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _810_
timestamp 1667941163
transform 1 0 19412 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _811_
timestamp 1667941163
transform 1 0 18584 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _812_
timestamp 1667941163
transform 1 0 18584 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _813_
timestamp 1667941163
transform 1 0 25668 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _814_
timestamp 1667941163
transform 1 0 24748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _815_
timestamp 1667941163
transform 1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _816_
timestamp 1667941163
transform 1 0 25760 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _817_
timestamp 1667941163
transform 1 0 25668 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _818_
timestamp 1667941163
transform 1 0 25668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _819_
timestamp 1667941163
transform 1 0 26128 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _820_
timestamp 1667941163
transform 1 0 25576 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _821_
timestamp 1667941163
transform 1 0 26128 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _822_
timestamp 1667941163
transform 1 0 25944 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _823_
timestamp 1667941163
transform 1 0 25300 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _824_
timestamp 1667941163
transform 1 0 26956 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _825_
timestamp 1667941163
transform 1 0 27140 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _826_
timestamp 1667941163
transform 1 0 27784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _827_
timestamp 1667941163
transform 1 0 29716 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _828_
timestamp 1667941163
transform 1 0 28980 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _829_
timestamp 1667941163
transform 1 0 28520 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _830_
timestamp 1667941163
transform 1 0 28796 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _831_
timestamp 1667941163
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _832_
timestamp 1667941163
transform 1 0 30820 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _833_
timestamp 1667941163
transform 1 0 30268 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _834_
timestamp 1667941163
transform 1 0 29900 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _835_
timestamp 1667941163
transform 1 0 24288 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _836_
timestamp 1667941163
transform 1 0 24840 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _837_
timestamp 1667941163
transform 1 0 25576 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _838_
timestamp 1667941163
transform 1 0 26312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _839_
timestamp 1667941163
transform 1 0 25760 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _840_
timestamp 1667941163
transform 1 0 25576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _841_
timestamp 1667941163
transform 1 0 23092 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _842_
timestamp 1667941163
transform 1 0 22632 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _843_
timestamp 1667941163
transform 1 0 23828 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _844_
timestamp 1667941163
transform 1 0 22264 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _845_
timestamp 1667941163
transform 1 0 22356 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _846_
timestamp 1667941163
transform 1 0 22172 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _847_
timestamp 1667941163
transform 1 0 21436 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _848_
timestamp 1667941163
transform 1 0 20516 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _849_
timestamp 1667941163
transform 1 0 20332 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _850_
timestamp 1667941163
transform 1 0 20608 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _851_
timestamp 1667941163
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _852_
timestamp 1667941163
transform 1 0 19688 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _853_
timestamp 1667941163
transform 1 0 20884 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _854_
timestamp 1667941163
transform 1 0 19964 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_1  _855_ pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 32844 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _856_
timestamp 1667941163
transform 1 0 31004 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _857_
timestamp 1667941163
transform 1 0 31372 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _858_
timestamp 1667941163
transform 1 0 32292 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _859_
timestamp 1667941163
transform 1 0 34868 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _860_
timestamp 1667941163
transform 1 0 35328 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _861_
timestamp 1667941163
transform 1 0 35512 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _862_
timestamp 1667941163
transform 1 0 36892 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _863_
timestamp 1667941163
transform 1 0 36892 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _864_
timestamp 1667941163
transform 1 0 32936 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _865_
timestamp 1667941163
transform 1 0 36708 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _866_
timestamp 1667941163
transform 1 0 34316 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _867_
timestamp 1667941163
transform 1 0 36616 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _868_
timestamp 1667941163
transform 1 0 36892 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _869_
timestamp 1667941163
transform 1 0 34868 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _870_
timestamp 1667941163
transform 1 0 36892 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _871_
timestamp 1667941163
transform 1 0 36892 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _872_
timestamp 1667941163
transform 1 0 36156 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _873_
timestamp 1667941163
transform 1 0 33396 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _874_
timestamp 1667941163
transform 1 0 35420 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _875_
timestamp 1667941163
transform 1 0 34868 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _876_
timestamp 1667941163
transform 1 0 35512 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _877_
timestamp 1667941163
transform 1 0 36708 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _878_
timestamp 1667941163
transform 1 0 36892 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _879_
timestamp 1667941163
transform 1 0 36892 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _880_
timestamp 1667941163
transform 1 0 35880 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _881_
timestamp 1667941163
transform 1 0 34868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _882_
timestamp 1667941163
transform 1 0 32292 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _883_
timestamp 1667941163
transform 1 0 31188 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _884_
timestamp 1667941163
transform 1 0 32016 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _885_
timestamp 1667941163
transform 1 0 30176 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _886_
timestamp 1667941163
transform 1 0 32016 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _887_
timestamp 1667941163
transform 1 0 34868 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _888_
timestamp 1667941163
transform 1 0 34868 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _889_
timestamp 1667941163
transform 1 0 34868 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _890_
timestamp 1667941163
transform 1 0 35236 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _891_
timestamp 1667941163
transform 1 0 27692 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _892_
timestamp 1667941163
transform 1 0 24196 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _893_
timestamp 1667941163
transform 1 0 25208 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _894_
timestamp 1667941163
transform 1 0 26404 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _895_
timestamp 1667941163
transform 1 0 28704 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _896_
timestamp 1667941163
transform 1 0 29716 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _897_
timestamp 1667941163
transform 1 0 28336 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _898_
timestamp 1667941163
transform 1 0 26404 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _899_
timestamp 1667941163
transform 1 0 27140 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _900_
timestamp 1667941163
transform 1 0 29992 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _901_
timestamp 1667941163
transform 1 0 22448 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _902_
timestamp 1667941163
transform 1 0 21988 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _903_
timestamp 1667941163
transform 1 0 22632 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _904_
timestamp 1667941163
transform 1 0 23460 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _905_
timestamp 1667941163
transform 1 0 22632 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _906_
timestamp 1667941163
transform 1 0 21712 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _907_
timestamp 1667941163
transform 1 0 22816 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _908_
timestamp 1667941163
transform 1 0 21436 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _909_
timestamp 1667941163
transform 1 0 34868 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _910_
timestamp 1667941163
transform 1 0 30176 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _911_
timestamp 1667941163
transform 1 0 32476 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _912_
timestamp 1667941163
transform 1 0 32660 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _913_
timestamp 1667941163
transform 1 0 30268 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _914_
timestamp 1667941163
transform 1 0 30176 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _915_
timestamp 1667941163
transform 1 0 30176 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _916_
timestamp 1667941163
transform 1 0 32016 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _917_
timestamp 1667941163
transform 1 0 32384 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _918_
timestamp 1667941163
transform 1 0 29624 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _919_
timestamp 1667941163
transform 1 0 30636 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _920_
timestamp 1667941163
transform 1 0 27784 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _921_
timestamp 1667941163
transform 1 0 26036 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _922_
timestamp 1667941163
transform 1 0 22080 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _923_
timestamp 1667941163
transform 1 0 23552 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _924_
timestamp 1667941163
transform 1 0 27140 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _925_
timestamp 1667941163
transform 1 0 29532 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _926_
timestamp 1667941163
transform 1 0 33580 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _927_
timestamp 1667941163
transform 1 0 32476 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _928_
timestamp 1667941163
transform 1 0 26496 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _929_
timestamp 1667941163
transform 1 0 28704 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _930_
timestamp 1667941163
transform 1 0 28796 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _931_
timestamp 1667941163
transform 1 0 24932 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _932_
timestamp 1667941163
transform 1 0 23920 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _933_
timestamp 1667941163
transform 1 0 22080 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _934_
timestamp 1667941163
transform 1 0 20056 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _935_
timestamp 1667941163
transform 1 0 19412 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _936_
timestamp 1667941163
transform 1 0 27600 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _937_
timestamp 1667941163
transform 1 0 31188 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _938_
timestamp 1667941163
transform 1 0 19780 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _939_
timestamp 1667941163
transform 1 0 19596 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _940_
timestamp 1667941163
transform 1 0 19872 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _941_
timestamp 1667941163
transform 1 0 19780 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _942_
timestamp 1667941163
transform 1 0 19688 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _943_
timestamp 1667941163
transform 1 0 19780 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _944_
timestamp 1667941163
transform 1 0 19780 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _945_
timestamp 1667941163
transform 1 0 19504 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _946_
timestamp 1667941163
transform 1 0 24288 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _947_
timestamp 1667941163
transform 1 0 23920 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _948_
timestamp 1667941163
transform 1 0 25024 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _949_
timestamp 1667941163
transform 1 0 25116 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _950_
timestamp 1667941163
transform 1 0 25300 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _951_
timestamp 1667941163
transform 1 0 27140 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _952_
timestamp 1667941163
transform 1 0 28980 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _953_
timestamp 1667941163
transform 1 0 29992 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _954_
timestamp 1667941163
transform 1 0 29808 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _955_
timestamp 1667941163
transform 1 0 24564 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _956_
timestamp 1667941163
transform 1 0 24564 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _957_
timestamp 1667941163
transform 1 0 23644 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _958_
timestamp 1667941163
transform 1 0 22540 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _959_
timestamp 1667941163
transform 1 0 21988 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _960_
timestamp 1667941163
transform 1 0 19872 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _961_
timestamp 1667941163
transform 1 0 19596 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _962_
timestamp 1667941163
transform 1 0 19504 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_1  _967_
timestamp 1667941163
transform 1 0 29900 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 29716 0 1 22848
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1667941163
transform 1 0 23368 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1667941163
transform 1 0 23368 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1667941163
transform 1 0 23368 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1667941163
transform 1 0 23368 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1667941163
transform 1 0 31188 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1667941163
transform 1 0 31188 0 1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1667941163
transform 1 0 31188 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1667941163
transform 1 0 33764 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1667941163
transform 1 0 1564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1667941163
transform 1 0 38088 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1667941163
transform 1 0 38088 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1667941163
transform 1 0 20056 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 1564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1667941163
transform 1 0 29716 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input7
timestamp 1667941163
transform 1 0 10396 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output8
timestamp 1667941163
transform 1 0 37996 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1667941163
transform 1 0 19412 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1667941163
transform 1 0 1564 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1667941163
transform 1 0 37996 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_12 pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1667941163
transform 1 0 9752 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_13
timestamp 1667941163
transform 1 0 29716 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_14
timestamp 1667941163
transform 1 0 1564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  rgb_mixer_15
timestamp 1667941163
transform 1 0 1564 0 1 20672
box -38 -48 314 592
<< labels >>
flabel metal3 s 39200 19048 39800 19168 0 FreeSans 480 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 662 39200 718 39800 0 FreeSans 224 90 0 0 enc0_a
port 1 nsew signal input
flabel metal3 s 39200 29248 39800 29368 0 FreeSans 480 0 0 0 enc0_b
port 2 nsew signal input
flabel metal2 s 38658 200 38714 800 0 FreeSans 224 90 0 0 enc1_a
port 3 nsew signal input
flabel metal2 s 19982 39200 20038 39800 0 FreeSans 224 90 0 0 enc1_b
port 4 nsew signal input
flabel metal2 s 18 200 74 800 0 FreeSans 224 90 0 0 enc2_a
port 5 nsew signal input
flabel metal2 s 28998 200 29054 800 0 FreeSans 224 90 0 0 enc2_b
port 6 nsew signal input
flabel metal2 s 9678 200 9734 800 0 FreeSans 224 90 0 0 io_oeb[0]
port 7 nsew signal tristate
flabel metal2 s 29642 39200 29698 39800 0 FreeSans 224 90 0 0 io_oeb[1]
port 8 nsew signal tristate
flabel metal3 s 200 10208 800 10328 0 FreeSans 480 0 0 0 io_oeb[2]
port 9 nsew signal tristate
flabel metal3 s 200 20408 800 20528 0 FreeSans 480 0 0 0 io_oeb[3]
port 10 nsew signal tristate
flabel metal2 s 39302 39200 39358 39800 0 FreeSans 224 90 0 0 pwm0_out
port 11 nsew signal tristate
flabel metal2 s 19338 200 19394 800 0 FreeSans 224 90 0 0 pwm1_out
port 12 nsew signal tristate
flabel metal3 s 200 30608 800 30728 0 FreeSans 480 0 0 0 pwm2_out
port 13 nsew signal tristate
flabel metal2 s 10322 39200 10378 39800 0 FreeSans 224 90 0 0 reset
port 14 nsew signal input
flabel metal3 s 39200 8848 39800 8968 0 FreeSans 480 0 0 0 sync
port 15 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 16 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 17 nsew ground bidirectional
rlabel metal1 19964 37536 19964 37536 0 vccd1
rlabel metal1 19964 36992 19964 36992 0 vssd1
rlabel metal2 33994 30498 33994 30498 0 _000_
rlabel via1 31321 30634 31321 30634 0 _001_
rlabel via1 31689 28526 31689 28526 0 _002_
rlabel metal1 32931 28118 32931 28118 0 _003_
rlabel metal2 34822 28322 34822 28322 0 _004_
rlabel via1 35645 30294 35645 30294 0 _005_
rlabel metal2 36754 31518 36754 31518 0 _006_
rlabel via1 37209 30702 37209 30702 0 _007_
rlabel metal1 37347 29614 37347 29614 0 _008_
rlabel metal2 34914 26044 34914 26044 0 _009_
rlabel metal2 36018 28322 36018 28322 0 _010_
rlabel metal1 35001 26962 35001 26962 0 _011_
rlabel metal1 36836 27438 36836 27438 0 _012_
rlabel metal1 36156 26010 36156 26010 0 _013_
rlabel metal1 34960 24922 34960 24922 0 _014_
rlabel metal1 37112 25262 37112 25262 0 _015_
rlabel metal2 37398 22610 37398 22610 0 _016_
rlabel metal2 36662 23970 36662 23970 0 _017_
rlabel metal1 34081 17238 34081 17238 0 _018_
rlabel metal1 35420 14586 35420 14586 0 _019_
rlabel metal2 34730 18734 34730 18734 0 _020_
rlabel via1 35829 19414 35829 19414 0 _021_
rlabel via1 37025 18734 37025 18734 0 _022_
rlabel metal1 37352 16966 37352 16966 0 _023_
rlabel metal2 38134 15266 38134 15266 0 _024_
rlabel metal1 36841 14382 36841 14382 0 _025_
rlabel metal1 35328 16966 35328 16966 0 _026_
rlabel via1 32609 22678 32609 22678 0 _027_
rlabel metal1 30252 27370 30252 27370 0 _028_
rlabel metal1 33258 24650 33258 24650 0 _029_
rlabel metal1 30953 23766 30953 23766 0 _030_
rlabel metal1 32236 24174 32236 24174 0 _031_
rlabel metal1 34990 23018 34990 23018 0 _032_
rlabel metal1 34714 22678 34714 22678 0 _033_
rlabel metal2 36018 20706 36018 20706 0 _034_
rlabel metal2 36662 21046 36662 21046 0 _035_
rlabel via1 28009 22610 28009 22610 0 _036_
rlabel metal1 25295 19414 25295 19414 0 _037_
rlabel via1 25525 20434 25525 20434 0 _038_
rlabel via1 26721 20842 26721 20842 0 _039_
rlabel metal1 28934 21998 28934 21998 0 _040_
rlabel metal1 29936 18258 29936 18258 0 _041_
rlabel metal1 28428 16762 28428 16762 0 _042_
rlabel metal1 28934 17850 28934 17850 0 _043_
rlabel metal1 27360 18258 27360 18258 0 _044_
rlabel metal1 32154 21896 32154 21896 0 _045_
rlabel metal1 23133 20842 23133 20842 0 _046_
rlabel metal1 22202 21590 22202 21590 0 _047_
rlabel via1 22949 23018 22949 23018 0 _048_
rlabel metal1 24564 24378 24564 24378 0 _049_
rlabel via1 22949 25262 22949 25262 0 _050_
rlabel metal2 22310 27642 22310 27642 0 _051_
rlabel metal1 22708 29206 22708 29206 0 _052_
rlabel via1 21753 30634 21753 30634 0 _053_
rlabel metal2 34638 29036 34638 29036 0 _054_
rlabel metal2 30038 14790 30038 14790 0 _055_
rlabel metal2 33442 19346 33442 19346 0 _056_
rlabel metal1 33069 20842 33069 20842 0 _057_
rlabel via1 30585 20910 30585 20910 0 _058_
rlabel via1 30493 17238 30493 17238 0 _059_
rlabel metal2 30590 16354 30590 16354 0 _060_
rlabel metal1 30820 15674 30820 15674 0 _061_
rlabel metal1 33391 18326 33391 18326 0 _062_
rlabel metal2 29762 31110 29762 31110 0 _063_
rlabel metal1 30856 31790 30856 31790 0 _064_
rlabel metal1 28060 32198 28060 32198 0 _065_
rlabel metal1 27135 31790 27135 31790 0 _066_
rlabel metal1 23501 31790 23501 31790 0 _067_
rlabel metal2 24978 30022 24978 30022 0 _068_
rlabel metal1 27094 29818 27094 29818 0 _069_
rlabel metal1 29752 29138 29752 29138 0 _070_
rlabel metal1 34403 14994 34403 14994 0 _071_
rlabel metal2 32430 31586 32430 31586 0 _072_
rlabel metal2 27186 16354 27186 16354 0 _073_
rlabel metal1 28658 15674 28658 15674 0 _074_
rlabel metal1 28842 13498 28842 13498 0 _075_
rlabel metal1 25208 14042 25208 14042 0 _076_
rlabel metal1 23736 14586 23736 14586 0 _077_
rlabel metal2 22954 14518 22954 14518 0 _078_
rlabel metal2 21298 14790 21298 14790 0 _079_
rlabel metal2 20470 14178 20470 14178 0 _080_
rlabel metal1 28658 20570 28658 20570 0 _081_
rlabel metal1 31086 14382 31086 14382 0 _082_
rlabel via1 20097 21522 20097 21522 0 _083_
rlabel metal1 19603 22678 19603 22678 0 _084_
rlabel metal1 19872 24378 19872 24378 0 _085_
rlabel via1 20097 25262 20097 25262 0 _086_
rlabel metal1 19304 27030 19304 27030 0 _087_
rlabel metal2 20194 28288 20194 28288 0 _088_
rlabel metal1 19504 29818 19504 29818 0 _089_
rlabel metal1 19734 30022 19734 30022 0 _090_
rlabel metal1 24702 22202 24702 22202 0 _091_
rlabel metal1 24467 27030 24467 27030 0 _092_
rlabel metal1 25525 28458 25525 28458 0 _093_
rlabel metal1 25525 26282 25525 26282 0 _094_
rlabel metal1 25520 24174 25520 24174 0 _095_
rlabel metal1 27687 24786 27687 24786 0 _096_
rlabel metal2 28566 24582 28566 24582 0 _097_
rlabel metal2 30866 24922 30866 24922 0 _098_
rlabel metal1 30171 25942 30171 25942 0 _099_
rlabel metal1 24656 20570 24656 20570 0 _100_
rlabel metal2 25622 18530 25622 18530 0 _101_
rlabel metal1 24789 16150 24789 16150 0 _102_
rlabel metal1 23179 18666 23179 18666 0 _103_
rlabel via1 22305 19414 22305 19414 0 _104_
rlabel metal2 20378 19618 20378 19618 0 _105_
rlabel metal1 19816 18734 19816 18734 0 _106_
rlabel metal1 19913 17238 19913 17238 0 _107_
rlabel metal1 33488 20434 33488 20434 0 _108_
rlabel metal1 33488 23086 33488 23086 0 _109_
rlabel metal1 30774 28662 30774 28662 0 _110_
rlabel via1 30408 28050 30408 28050 0 _111_
rlabel metal1 32085 25942 32085 25942 0 _112_
rlabel metal1 28957 26962 28957 26962 0 _113_
rlabel metal1 28198 27030 28198 27030 0 _114_
rlabel metal2 27738 26996 27738 26996 0 _115_
rlabel metal1 27370 27098 27370 27098 0 _116_
rlabel metal1 28014 29104 28014 29104 0 _117_
rlabel metal1 27646 28458 27646 28458 0 _118_
rlabel metal1 27186 28186 27186 28186 0 _119_
rlabel metal2 28014 28220 28014 28220 0 _120_
rlabel metal1 28382 28186 28382 28186 0 _121_
rlabel metal1 27186 27642 27186 27642 0 _122_
rlabel metal2 27554 27914 27554 27914 0 _123_
rlabel metal2 28198 27132 28198 27132 0 _124_
rlabel metal1 29302 27098 29302 27098 0 _125_
rlabel metal2 30498 27778 30498 27778 0 _126_
rlabel metal1 30636 28186 30636 28186 0 _127_
rlabel metal2 32522 36317 32522 36317 0 _128_
rlabel metal1 20194 16218 20194 16218 0 _129_
rlabel metal1 21114 16048 21114 16048 0 _130_
rlabel metal2 20930 15878 20930 15878 0 _131_
rlabel metal2 23506 16592 23506 16592 0 _132_
rlabel metal1 24426 15402 24426 15402 0 _133_
rlabel metal2 23138 16082 23138 16082 0 _134_
rlabel metal2 25530 15844 25530 15844 0 _135_
rlabel metal1 25254 16524 25254 16524 0 _136_
rlabel metal1 26082 16116 26082 16116 0 _137_
rlabel metal1 25254 16218 25254 16218 0 _138_
rlabel metal1 25162 16762 25162 16762 0 _139_
rlabel metal1 23368 16558 23368 16558 0 _140_
rlabel metal1 22034 16490 22034 16490 0 _141_
rlabel metal1 20746 16150 20746 16150 0 _142_
rlabel metal1 21390 15912 21390 15912 0 _143_
rlabel metal1 20470 15946 20470 15946 0 _144_
rlabel metal1 20056 20230 20056 20230 0 _145_
rlabel metal2 20378 30192 20378 30192 0 _146_
rlabel metal1 21620 29682 21620 29682 0 _147_
rlabel metal2 21850 28458 21850 28458 0 _148_
rlabel metal2 21390 26690 21390 26690 0 _149_
rlabel metal1 22586 24854 22586 24854 0 _150_
rlabel metal1 22126 24718 22126 24718 0 _151_
rlabel metal1 21759 24208 21759 24208 0 _152_
rlabel metal2 21666 23290 21666 23290 0 _153_
rlabel via1 21947 23086 21947 23086 0 _154_
rlabel metal1 21712 23290 21712 23290 0 _155_
rlabel metal2 21666 24004 21666 24004 0 _156_
rlabel metal1 21666 25296 21666 25296 0 _157_
rlabel metal1 22034 26928 22034 26928 0 _158_
rlabel metal1 21666 28594 21666 28594 0 _159_
rlabel metal1 21758 29546 21758 29546 0 _160_
rlabel metal1 22356 29818 22356 29818 0 _161_
rlabel metal1 34835 18258 34835 18258 0 _162_
rlabel metal1 36570 30090 36570 30090 0 _163_
rlabel metal1 34270 29818 34270 29818 0 _164_
rlabel metal2 34270 29410 34270 29410 0 _165_
rlabel metal1 36179 29478 36179 29478 0 _166_
rlabel metal1 35052 29818 35052 29818 0 _167_
rlabel metal2 34362 27846 34362 27846 0 _168_
rlabel metal1 22862 32198 22862 32198 0 _169_
rlabel metal1 26680 31994 26680 31994 0 _170_
rlabel metal2 31786 29308 31786 29308 0 _171_
rlabel metal1 37674 25806 37674 25806 0 _172_
rlabel metal2 33442 28764 33442 28764 0 _173_
rlabel metal2 35006 28220 35006 28220 0 _174_
rlabel metal1 35696 29274 35696 29274 0 _175_
rlabel metal1 36662 30906 36662 30906 0 _176_
rlabel metal1 37766 31450 37766 31450 0 _177_
rlabel metal2 37858 30532 37858 30532 0 _178_
rlabel metal1 34500 27098 34500 27098 0 _179_
rlabel metal1 37674 24650 37674 24650 0 _180_
rlabel metal1 35098 26418 35098 26418 0 _181_
rlabel metal2 36478 27132 36478 27132 0 _182_
rlabel metal1 36754 26826 36754 26826 0 _183_
rlabel metal2 36202 26588 36202 26588 0 _184_
rlabel metal2 36202 28492 36202 28492 0 _185_
rlabel metal1 37720 27098 37720 27098 0 _186_
rlabel metal1 36892 26010 36892 26010 0 _187_
rlabel metal1 35236 24786 35236 24786 0 _188_
rlabel metal1 36938 25908 36938 25908 0 _189_
rlabel metal2 37674 22100 37674 22100 0 _190_
rlabel metal2 37582 22746 37582 22746 0 _191_
rlabel metal1 37582 22746 37582 22746 0 _192_
rlabel metal2 34730 19516 34730 19516 0 _193_
rlabel metal1 37636 18326 37636 18326 0 _194_
rlabel metal1 34638 18190 34638 18190 0 _195_
rlabel metal2 36846 17918 36846 17918 0 _196_
rlabel metal2 35558 17476 35558 17476 0 _197_
rlabel metal1 35328 17850 35328 17850 0 _198_
rlabel metal2 35466 14212 35466 14212 0 _199_
rlabel metal2 36018 19108 36018 19108 0 _200_
rlabel metal1 37306 17850 37306 17850 0 _201_
rlabel metal2 37674 17340 37674 17340 0 _202_
rlabel metal2 38318 15436 38318 15436 0 _203_
rlabel metal2 37674 15164 37674 15164 0 _204_
rlabel metal1 35650 16218 35650 16218 0 _205_
rlabel metal1 33764 26282 33764 26282 0 _206_
rlabel metal2 35558 22508 35558 22508 0 _207_
rlabel metal2 34270 23426 34270 23426 0 _208_
rlabel metal2 33074 23834 33074 23834 0 _209_
rlabel metal2 35650 22134 35650 22134 0 _210_
rlabel metal1 32844 23222 32844 23222 0 _211_
rlabel metal2 29210 27676 29210 27676 0 _212_
rlabel metal2 31786 22950 31786 22950 0 _213_
rlabel metal1 31280 24174 31280 24174 0 _214_
rlabel metal2 32338 24004 32338 24004 0 _215_
rlabel metal1 34684 24174 34684 24174 0 _216_
rlabel metal1 34408 22202 34408 22202 0 _217_
rlabel metal2 36202 20876 36202 20876 0 _218_
rlabel metal1 36846 20468 36846 20468 0 _219_
rlabel metal2 20102 29410 20102 29410 0 _220_
rlabel metal2 28842 20230 28842 20230 0 _221_
rlabel metal1 28520 21114 28520 21114 0 _222_
rlabel metal1 28474 19482 28474 19482 0 _223_
rlabel metal2 28658 20162 28658 20162 0 _224_
rlabel metal1 30866 21998 30866 21998 0 _225_
rlabel metal1 28106 20230 28106 20230 0 _226_
rlabel metal1 24426 15878 24426 15878 0 _227_
rlabel metal2 26266 20774 26266 20774 0 _228_
rlabel metal1 26634 21556 26634 21556 0 _229_
rlabel metal1 28980 21658 28980 21658 0 _230_
rlabel metal2 29486 19516 29486 19516 0 _231_
rlabel metal1 33626 17612 33626 17612 0 _232_
rlabel metal1 28750 16558 28750 16558 0 _233_
rlabel metal1 29946 17612 29946 17612 0 _234_
rlabel metal1 27186 17850 27186 17850 0 _235_
rlabel metal1 33948 20434 33948 20434 0 _236_
rlabel metal2 32890 18394 32890 18394 0 _237_
rlabel metal2 33626 20740 33626 20740 0 _238_
rlabel metal1 32706 20570 32706 20570 0 _239_
rlabel metal1 32752 19482 32752 19482 0 _240_
rlabel metal1 32476 21658 32476 21658 0 _241_
rlabel metal1 20976 21930 20976 21930 0 _242_
rlabel metal1 22310 22032 22310 22032 0 _243_
rlabel metal1 23644 22610 23644 22610 0 _244_
rlabel metal2 23138 24684 23138 24684 0 _245_
rlabel metal2 24794 24684 24794 24684 0 _246_
rlabel metal2 24610 24786 24610 24786 0 _247_
rlabel metal2 23138 26180 23138 26180 0 _248_
rlabel metal1 25024 25466 25024 25466 0 _249_
rlabel metal1 23644 28186 23644 28186 0 _250_
rlabel metal2 23598 27778 23598 27778 0 _251_
rlabel metal2 22402 30124 22402 30124 0 _252_
rlabel metal2 23782 29002 23782 29002 0 _253_
rlabel metal1 22586 31314 22586 31314 0 _254_
rlabel metal1 30176 13498 30176 13498 0 _255_
rlabel metal1 33396 18734 33396 18734 0 _256_
rlabel metal1 31234 20570 31234 20570 0 _257_
rlabel metal2 30958 19516 30958 19516 0 _258_
rlabel metal2 30774 16796 30774 16796 0 _259_
rlabel metal2 30958 15674 30958 15674 0 _260_
rlabel metal1 34040 17850 34040 17850 0 _261_
rlabel metal1 34730 32946 34730 32946 0 _262_
rlabel metal2 33994 33184 33994 33184 0 _263_
rlabel metal1 34362 32266 34362 32266 0 _264_
rlabel metal1 33626 32470 33626 32470 0 _265_
rlabel metal1 32522 32946 32522 32946 0 _266_
rlabel metal1 25484 31858 25484 31858 0 _267_
rlabel metal1 29946 30736 29946 30736 0 _268_
rlabel metal2 30406 32674 30406 32674 0 _269_
rlabel metal2 30590 33660 30590 33660 0 _270_
rlabel metal1 30360 33966 30360 33966 0 _271_
rlabel metal2 31234 33490 31234 33490 0 _272_
rlabel metal1 31372 33082 31372 33082 0 _273_
rlabel metal1 30820 32402 30820 32402 0 _274_
rlabel metal2 25254 32028 25254 32028 0 _275_
rlabel metal1 28474 33490 28474 33490 0 _276_
rlabel metal2 29210 33524 29210 33524 0 _277_
rlabel metal1 26082 32334 26082 32334 0 _278_
rlabel metal1 28198 34034 28198 34034 0 _279_
rlabel metal2 28474 33626 28474 33626 0 _280_
rlabel metal2 29118 32878 29118 32878 0 _281_
rlabel metal1 28474 32368 28474 32368 0 _282_
rlabel metal2 26542 33796 26542 33796 0 _283_
rlabel metal1 27232 34102 27232 34102 0 _284_
rlabel metal1 26772 33082 26772 33082 0 _285_
rlabel metal2 28382 32810 28382 32810 0 _286_
rlabel metal1 27692 33082 27692 33082 0 _287_
rlabel metal2 25162 33116 25162 33116 0 _288_
rlabel metal2 24886 33252 24886 33252 0 _289_
rlabel metal1 23046 32946 23046 32946 0 _290_
rlabel metal1 23828 32878 23828 32878 0 _291_
rlabel metal2 25070 32300 25070 32300 0 _292_
rlabel metal2 25254 32708 25254 32708 0 _293_
rlabel metal2 23782 32674 23782 32674 0 _294_
rlabel metal1 24426 29614 24426 29614 0 _295_
rlabel metal2 24886 30192 24886 30192 0 _296_
rlabel metal1 25530 30668 25530 30668 0 _297_
rlabel metal2 25806 30192 25806 30192 0 _298_
rlabel metal2 26082 30022 26082 30022 0 _299_
rlabel metal2 25990 32708 25990 32708 0 _300_
rlabel metal1 25300 30906 25300 30906 0 _301_
rlabel metal1 26450 30090 26450 30090 0 _302_
rlabel metal1 27232 29614 27232 29614 0 _303_
rlabel metal2 29394 30532 29394 30532 0 _304_
rlabel metal2 29486 29682 29486 29682 0 _305_
rlabel metal1 28796 29274 28796 29274 0 _306_
rlabel metal2 28750 29852 28750 29852 0 _307_
rlabel metal1 34638 15470 34638 15470 0 _308_
rlabel metal1 32614 31348 32614 31348 0 _309_
rlabel metal1 33810 16082 33810 16082 0 _310_
rlabel metal1 32982 16150 32982 16150 0 _311_
rlabel metal1 32982 15504 32982 15504 0 _312_
rlabel metal2 33028 15470 33028 15470 0 _313_
rlabel metal2 21206 14654 21206 14654 0 _314_
rlabel metal1 25530 13974 25530 13974 0 _315_
rlabel metal2 27370 16524 27370 16524 0 _316_
rlabel metal2 32706 15334 32706 15334 0 _317_
rlabel metal1 27646 15028 27646 15028 0 _318_
rlabel metal2 27738 15300 27738 15300 0 _319_
rlabel metal1 26726 15538 26726 15538 0 _320_
rlabel metal2 27830 15130 27830 15130 0 _321_
rlabel metal1 27002 15436 27002 15436 0 _322_
rlabel metal1 26174 12172 26174 12172 0 _323_
rlabel metal2 28382 13260 28382 13260 0 _324_
rlabel metal1 19596 12206 19596 12206 0 _325_
rlabel via1 27370 12415 27370 12415 0 _326_
rlabel metal2 26818 12784 26818 12784 0 _327_
rlabel metal2 28014 13906 28014 13906 0 _328_
rlabel metal2 29026 13838 29026 13838 0 _329_
rlabel metal1 26312 12342 26312 12342 0 _330_
rlabel metal1 26082 13260 26082 13260 0 _331_
rlabel metal1 25484 13362 25484 13362 0 _332_
rlabel metal1 25300 13498 25300 13498 0 _333_
rlabel metal2 26450 12410 26450 12410 0 _334_
rlabel metal2 24794 12614 24794 12614 0 _335_
rlabel metal1 23690 12342 23690 12342 0 _336_
rlabel metal1 23966 12954 23966 12954 0 _337_
rlabel metal1 23690 13260 23690 13260 0 _338_
rlabel metal1 24104 14042 24104 14042 0 _339_
rlabel metal1 22586 12308 22586 12308 0 _340_
rlabel metal1 23184 13294 23184 13294 0 _341_
rlabel metal2 22402 13430 22402 13430 0 _342_
rlabel metal1 22770 13498 22770 13498 0 _343_
rlabel metal1 20976 12410 20976 12410 0 _344_
rlabel metal1 20056 12410 20056 12410 0 _345_
rlabel metal2 20838 12036 20838 12036 0 _346_
rlabel metal1 23322 12614 23322 12614 0 _347_
rlabel metal1 20976 12274 20976 12274 0 _348_
rlabel metal1 21068 13294 21068 13294 0 _349_
rlabel metal2 21298 13872 21298 13872 0 _350_
rlabel metal1 20424 12954 20424 12954 0 _351_
rlabel metal1 19734 13702 19734 13702 0 _352_
rlabel metal1 19964 13498 19964 13498 0 _353_
rlabel metal1 20010 13872 20010 13872 0 _354_
rlabel metal1 30314 15504 30314 15504 0 _355_
rlabel metal1 26680 23698 26680 23698 0 _356_
rlabel metal2 26358 22950 26358 22950 0 _357_
rlabel metal1 26082 23120 26082 23120 0 _358_
rlabel metal1 26174 23052 26174 23052 0 _359_
rlabel metal1 21344 21998 21344 21998 0 _360_
rlabel metal1 19136 29138 19136 29138 0 _361_
rlabel metal1 20286 22032 20286 22032 0 _362_
rlabel metal1 19642 23766 19642 23766 0 _363_
rlabel metal1 18722 22202 18722 22202 0 _364_
rlabel metal1 18262 21998 18262 21998 0 _365_
rlabel metal1 18262 21522 18262 21522 0 _366_
rlabel metal1 18860 21862 18860 21862 0 _367_
rlabel metal1 18998 21658 18998 21658 0 _368_
rlabel metal2 17894 23460 17894 23460 0 _369_
rlabel metal1 18860 24174 18860 24174 0 _370_
rlabel metal2 17250 24038 17250 24038 0 _371_
rlabel metal1 18032 24718 18032 24718 0 _372_
rlabel metal1 17986 24276 17986 24276 0 _373_
rlabel metal1 18768 23698 18768 23698 0 _374_
rlabel metal1 19734 23834 19734 23834 0 _375_
rlabel metal1 18860 25330 18860 25330 0 _376_
rlabel metal1 18860 24786 18860 24786 0 _377_
rlabel metal2 18630 24956 18630 24956 0 _378_
rlabel metal1 19136 24650 19136 24650 0 _379_
rlabel metal1 17434 24378 17434 24378 0 _380_
rlabel metal1 18078 26316 18078 26316 0 _381_
rlabel metal1 17250 27506 17250 27506 0 _382_
rlabel metal2 18538 26554 18538 26554 0 _383_
rlabel metal1 18492 26554 18492 26554 0 _384_
rlabel metal1 18906 26554 18906 26554 0 _385_
rlabel metal1 17526 27982 17526 27982 0 _386_
rlabel metal2 18446 27812 18446 27812 0 _387_
rlabel metal1 19320 27914 19320 27914 0 _388_
rlabel metal1 20332 27914 20332 27914 0 _389_
rlabel metal1 17204 30022 17204 30022 0 _390_
rlabel metal1 16790 29818 16790 29818 0 _391_
rlabel metal2 17250 30090 17250 30090 0 _392_
rlabel metal1 17572 27098 17572 27098 0 _393_
rlabel metal2 17342 28288 17342 28288 0 _394_
rlabel metal2 18722 29308 18722 29308 0 _395_
rlabel metal1 19550 29274 19550 29274 0 _396_
rlabel metal2 18630 29444 18630 29444 0 _397_
rlabel metal1 19458 29750 19458 29750 0 _398_
rlabel metal1 18814 30260 18814 30260 0 _399_
rlabel metal1 18860 29818 18860 29818 0 _400_
rlabel metal1 24978 22032 24978 22032 0 _401_
rlabel metal2 25806 28662 25806 28662 0 _402_
rlabel metal2 25714 26724 25714 26724 0 _403_
rlabel metal1 26450 25262 26450 25262 0 _404_
rlabel metal2 26542 24752 26542 24752 0 _405_
rlabel metal1 25346 24718 25346 24718 0 _406_
rlabel metal1 28014 25296 28014 25296 0 _407_
rlabel metal1 27600 24378 27600 24378 0 _408_
rlabel metal1 29026 23732 29026 23732 0 _409_
rlabel metal1 28934 23834 28934 23834 0 _410_
rlabel metal1 29624 25126 29624 25126 0 _411_
rlabel metal1 30820 24786 30820 24786 0 _412_
rlabel metal2 30130 26554 30130 26554 0 _413_
rlabel metal2 25806 19108 25806 19108 0 _414_
rlabel metal1 26036 17034 26036 17034 0 _415_
rlabel metal1 25898 17170 25898 17170 0 _416_
rlabel metal1 23782 17850 23782 17850 0 _417_
rlabel metal1 23414 17306 23414 17306 0 _418_
rlabel metal2 21666 19244 21666 19244 0 _419_
rlabel metal1 22448 18394 22448 18394 0 _420_
rlabel metal1 20930 18666 20930 18666 0 _421_
rlabel metal2 20562 19788 20562 19788 0 _422_
rlabel metal1 20562 17850 20562 17850 0 _423_
rlabel metal2 20194 18836 20194 18836 0 _424_
rlabel metal1 20194 17680 20194 17680 0 _425_
rlabel metal3 37567 19108 37567 19108 0 clk
rlabel metal2 33810 23494 33810 23494 0 clknet_0_clk
rlabel metal1 19550 18734 19550 18734 0 clknet_3_0__leaf_clk
rlabel metal1 27094 20910 27094 20910 0 clknet_3_1__leaf_clk
rlabel metal1 21758 31858 21758 31858 0 clknet_3_2__leaf_clk
rlabel metal1 26128 28526 26128 28526 0 clknet_3_3__leaf_clk
rlabel metal1 32062 16694 32062 16694 0 clknet_3_4__leaf_clk
rlabel metal1 36938 16694 36938 16694 0 clknet_3_5__leaf_clk
rlabel metal2 32522 31246 32522 31246 0 clknet_3_6__leaf_clk
rlabel metal1 36846 25330 36846 25330 0 clknet_3_7__leaf_clk
rlabel metal2 31878 30090 31878 30090 0 debounce0_a.button_hist\[0\]
rlabel metal2 32798 28934 32798 28934 0 debounce0_a.button_hist\[1\]
rlabel metal1 33994 29206 33994 29206 0 debounce0_a.button_hist\[2\]
rlabel metal2 35374 28764 35374 28764 0 debounce0_a.button_hist\[3\]
rlabel metal1 36754 30328 36754 30328 0 debounce0_a.button_hist\[4\]
rlabel metal1 37444 30090 37444 30090 0 debounce0_a.button_hist\[5\]
rlabel metal1 37904 30362 37904 30362 0 debounce0_a.button_hist\[6\]
rlabel metal1 37628 29818 37628 29818 0 debounce0_a.button_hist\[7\]
rlabel metal1 34178 30566 34178 30566 0 debounce0_a.debounced
rlabel metal1 35604 27642 35604 27642 0 debounce0_b.button_hist\[0\]
rlabel metal1 37490 27030 37490 27030 0 debounce0_b.button_hist\[1\]
rlabel metal2 36386 26758 36386 26758 0 debounce0_b.button_hist\[2\]
rlabel metal1 38318 26418 38318 26418 0 debounce0_b.button_hist\[3\]
rlabel metal1 37444 24922 37444 24922 0 debounce0_b.button_hist\[4\]
rlabel metal1 37214 24786 37214 24786 0 debounce0_b.button_hist\[5\]
rlabel metal1 37260 24854 37260 24854 0 debounce0_b.button_hist\[6\]
rlabel metal1 37766 24752 37766 24752 0 debounce0_b.button_hist\[7\]
rlabel metal2 36662 26384 36662 26384 0 debounce0_b.debounced
rlabel metal2 36570 17765 36570 17765 0 debounce1_a.button_hist\[0\]
rlabel metal1 36662 18292 36662 18292 0 debounce1_a.button_hist\[1\]
rlabel metal2 36662 18394 36662 18394 0 debounce1_a.button_hist\[2\]
rlabel metal2 37490 18122 37490 18122 0 debounce1_a.button_hist\[3\]
rlabel metal1 37490 16116 37490 16116 0 debounce1_a.button_hist\[4\]
rlabel metal1 36524 17034 36524 17034 0 debounce1_a.button_hist\[5\]
rlabel metal1 36846 17238 36846 17238 0 debounce1_a.button_hist\[6\]
rlabel metal2 36294 16898 36294 16898 0 debounce1_a.button_hist\[7\]
rlabel metal2 34822 17442 34822 17442 0 debounce1_a.debounced
rlabel metal1 33028 26418 33028 26418 0 debounce1_b.button_hist\[0\]
rlabel metal1 33672 25126 33672 25126 0 debounce1_b.button_hist\[1\]
rlabel metal1 33028 23154 33028 23154 0 debounce1_b.button_hist\[2\]
rlabel metal2 33442 24548 33442 24548 0 debounce1_b.button_hist\[3\]
rlabel metal1 34638 21930 34638 21930 0 debounce1_b.button_hist\[4\]
rlabel metal2 36294 22202 36294 22202 0 debounce1_b.button_hist\[5\]
rlabel metal2 35282 20604 35282 20604 0 debounce1_b.button_hist\[6\]
rlabel metal2 36202 21862 36202 21862 0 debounce1_b.button_hist\[7\]
rlabel metal2 33718 22882 33718 22882 0 debounce1_b.debounced
rlabel metal2 28014 20604 28014 20604 0 debounce2_a.button_hist\[0\]
rlabel metal1 27278 20434 27278 20434 0 debounce2_a.button_hist\[1\]
rlabel metal2 28658 21182 28658 21182 0 debounce2_a.button_hist\[2\]
rlabel metal1 28520 19822 28520 19822 0 debounce2_a.button_hist\[3\]
rlabel metal2 28842 18020 28842 18020 0 debounce2_a.button_hist\[4\]
rlabel metal2 28290 18020 28290 18020 0 debounce2_a.button_hist\[5\]
rlabel metal1 27784 18598 27784 18598 0 debounce2_a.button_hist\[6\]
rlabel metal1 28474 18734 28474 18734 0 debounce2_a.button_hist\[7\]
rlabel metal1 29118 22508 29118 22508 0 debounce2_a.debounced
rlabel metal2 33258 19465 33258 19465 0 debounce2_b.button_hist\[0\]
rlabel metal2 33258 20196 33258 20196 0 debounce2_b.button_hist\[1\]
rlabel metal2 32522 21250 32522 21250 0 debounce2_b.button_hist\[2\]
rlabel metal1 32522 20332 32522 20332 0 debounce2_b.button_hist\[3\]
rlabel metal2 32522 18190 32522 18190 0 debounce2_b.button_hist\[4\]
rlabel metal1 32338 17272 32338 17272 0 debounce2_b.button_hist\[5\]
rlabel metal1 32706 17136 32706 17136 0 debounce2_b.button_hist\[6\]
rlabel metal1 32614 17204 32614 17204 0 debounce2_b.button_hist\[7\]
rlabel metal1 32798 21556 32798 21556 0 debounce2_b.debounced
rlabel metal1 1242 37230 1242 37230 0 enc0_a
rlabel metal2 38318 30549 38318 30549 0 enc0_b
rlabel metal2 38686 1588 38686 1588 0 enc1_a
rlabel metal1 20148 37230 20148 37230 0 enc1_b
rlabel metal2 46 1588 46 1588 0 enc2_a
rlabel metal2 29026 1588 29026 1588 0 enc2_b
rlabel metal2 36294 32164 36294 32164 0 encoder0.old_a
rlabel metal2 34454 32164 34454 32164 0 encoder0.old_b
rlabel metal1 30360 33490 30360 33490 0 encoder0.value\[0\]
rlabel metal1 30360 32402 30360 32402 0 encoder0.value\[1\]
rlabel metal1 28290 32470 28290 32470 0 encoder0.value\[2\]
rlabel metal1 27416 32878 27416 32878 0 encoder0.value\[3\]
rlabel metal1 24012 32742 24012 32742 0 encoder0.value\[4\]
rlabel metal1 25438 32402 25438 32402 0 encoder0.value\[5\]
rlabel via1 30038 28050 30038 28050 0 encoder0.value\[6\]
rlabel metal1 29486 29614 29486 29614 0 encoder0.value\[7\]
rlabel metal1 33258 14994 33258 14994 0 encoder1.old_a
rlabel metal2 32614 14756 32614 14756 0 encoder1.old_b
rlabel metal1 27922 16456 27922 16456 0 encoder1.value\[0\]
rlabel metal1 29256 14994 29256 14994 0 encoder1.value\[1\]
rlabel via1 26358 12699 26358 12699 0 encoder1.value\[2\]
rlabel metal1 25852 12818 25852 12818 0 encoder1.value\[3\]
rlabel metal1 24472 15470 24472 15470 0 encoder1.value\[4\]
rlabel metal1 22494 12206 22494 12206 0 encoder1.value\[5\]
rlabel metal1 21528 12206 21528 12206 0 encoder1.value\[6\]
rlabel metal1 20654 13294 20654 13294 0 encoder1.value\[7\]
rlabel metal1 26910 23188 26910 23188 0 encoder2.old_a
rlabel metal2 25714 22848 25714 22848 0 encoder2.old_b
rlabel metal1 18446 21896 18446 21896 0 encoder2.value\[0\]
rlabel metal1 21160 22746 21160 22746 0 encoder2.value\[1\]
rlabel metal1 16698 24378 16698 24378 0 encoder2.value\[2\]
rlabel metal1 17296 25874 17296 25874 0 encoder2.value\[3\]
rlabel metal2 21114 26554 21114 26554 0 encoder2.value\[4\]
rlabel metal2 17158 27506 17158 27506 0 encoder2.value\[5\]
rlabel metal2 17158 29954 17158 29954 0 encoder2.value\[6\]
rlabel metal2 20286 30906 20286 30906 0 encoder2.value\[7\]
rlabel metal2 1610 34442 1610 34442 0 net1
rlabel metal2 1610 30124 1610 30124 0 net10
rlabel metal1 33994 8942 33994 8942 0 net11
rlabel metal2 9706 1588 9706 1588 0 net12
rlabel metal1 29808 37434 29808 37434 0 net13
rlabel metal3 1234 10268 1234 10268 0 net14
rlabel metal3 1234 20468 1234 20468 0 net15
rlabel metal1 36938 29138 36938 29138 0 net2
rlabel metal1 37076 13906 37076 13906 0 net3
rlabel metal1 22310 37094 22310 37094 0 net4
rlabel metal2 1886 9078 1886 9078 0 net5
rlabel metal1 29716 2618 29716 2618 0 net6
rlabel metal2 10626 32640 10626 32640 0 net7
rlabel metal2 32338 37060 32338 37060 0 net8
rlabel metal2 19458 4657 19458 4657 0 net9
rlabel metal1 26726 28050 26726 28050 0 pwm0.count\[0\]
rlabel metal2 26450 28934 26450 28934 0 pwm0.count\[1\]
rlabel metal2 26174 27200 26174 27200 0 pwm0.count\[2\]
rlabel metal2 27186 25908 27186 25908 0 pwm0.count\[3\]
rlabel metal2 28566 25636 28566 25636 0 pwm0.count\[4\]
rlabel metal2 29026 25908 29026 25908 0 pwm0.count\[5\]
rlabel metal2 31418 25670 31418 25670 0 pwm0.count\[6\]
rlabel metal2 31050 28288 31050 28288 0 pwm0.count\[7\]
rlabel metal1 38778 37434 38778 37434 0 pwm0_out
rlabel metal2 25162 20094 25162 20094 0 pwm1.count\[0\]
rlabel metal2 25990 19312 25990 19312 0 pwm1.count\[1\]
rlabel metal2 25346 16252 25346 16252 0 pwm1.count\[2\]
rlabel metal2 22678 16320 22678 16320 0 pwm1.count\[3\]
rlabel metal2 22402 18700 22402 18700 0 pwm1.count\[4\]
rlabel metal1 21160 16150 21160 16150 0 pwm1.count\[5\]
rlabel metal1 20470 16524 20470 16524 0 pwm1.count\[6\]
rlabel metal1 20562 16966 20562 16966 0 pwm1.count\[7\]
rlabel metal2 19366 1520 19366 1520 0 pwm1_out
rlabel metal1 23200 22678 23200 22678 0 pwm2.count\[0\]
rlabel metal1 21574 23052 21574 23052 0 pwm2.count\[1\]
rlabel metal1 21942 24072 21942 24072 0 pwm2.count\[2\]
rlabel metal1 24702 24922 24702 24922 0 pwm2.count\[3\]
rlabel metal1 24058 25364 24058 25364 0 pwm2.count\[4\]
rlabel metal1 22816 28730 22816 28730 0 pwm2.count\[5\]
rlabel metal1 22011 29614 22011 29614 0 pwm2.count\[6\]
rlabel metal2 22862 31076 22862 31076 0 pwm2.count\[7\]
rlabel metal3 1234 30668 1234 30668 0 pwm2_out
rlabel metal1 10442 37230 10442 37230 0 reset
rlabel metal2 38226 8857 38226 8857 0 sync
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
