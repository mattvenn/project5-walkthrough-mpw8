magic
tech sky130A
magscale 1 2
timestamp 1672748043
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 39362 37584
<< metal2 >>
rect 662 39200 718 39800
rect 10322 39200 10378 39800
rect 19982 39200 20038 39800
rect 29642 39200 29698 39800
rect 39302 39200 39358 39800
rect 18 200 74 800
rect 9678 200 9734 800
rect 19338 200 19394 800
rect 28998 200 29054 800
rect 38658 200 38714 800
<< obsm2 >>
rect 20 39144 606 39200
rect 774 39144 10266 39200
rect 10434 39144 19926 39200
rect 20094 39144 29586 39200
rect 29754 39144 39246 39200
rect 20 856 39356 39144
rect 130 800 9622 856
rect 9790 800 19282 856
rect 19450 800 28942 856
rect 29110 800 38602 856
rect 38770 800 39356 856
<< metal3 >>
rect 200 30608 800 30728
rect 39200 29248 39800 29368
rect 200 20408 800 20528
rect 39200 19048 39800 19168
rect 200 10208 800 10328
rect 39200 8848 39800 8968
<< obsm3 >>
rect 800 30808 39200 37569
rect 880 30528 39200 30808
rect 800 29448 39200 30528
rect 800 29168 39120 29448
rect 800 20608 39200 29168
rect 880 20328 39200 20608
rect 800 19248 39200 20328
rect 800 18968 39120 19248
rect 800 10408 39200 18968
rect 880 10128 39200 10408
rect 800 9048 39200 10128
rect 800 8768 39120 9048
rect 800 2143 39200 8768
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal3 s 39200 19048 39800 19168 6 clk
port 1 nsew signal input
rlabel metal2 s 662 39200 718 39800 6 enc0_a
port 2 nsew signal input
rlabel metal3 s 39200 29248 39800 29368 6 enc0_b
port 3 nsew signal input
rlabel metal2 s 38658 200 38714 800 6 enc1_a
port 4 nsew signal input
rlabel metal2 s 19982 39200 20038 39800 6 enc1_b
port 5 nsew signal input
rlabel metal2 s 18 200 74 800 6 enc2_a
port 6 nsew signal input
rlabel metal2 s 28998 200 29054 800 6 enc2_b
port 7 nsew signal input
rlabel metal2 s 9678 200 9734 800 6 io_oeb[0]
port 8 nsew signal output
rlabel metal2 s 29642 39200 29698 39800 6 io_oeb[1]
port 9 nsew signal output
rlabel metal3 s 200 10208 800 10328 6 io_oeb[2]
port 10 nsew signal output
rlabel metal3 s 200 20408 800 20528 6 io_oeb[3]
port 11 nsew signal output
rlabel metal2 s 39302 39200 39358 39800 6 pwm0_out
port 12 nsew signal output
rlabel metal2 s 19338 200 19394 800 6 pwm1_out
port 13 nsew signal output
rlabel metal3 s 200 30608 800 30728 6 pwm2_out
port 14 nsew signal output
rlabel metal2 s 10322 39200 10378 39800 6 reset
port 15 nsew signal input
rlabel metal3 s 39200 8848 39800 8968 6 sync
port 16 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 17 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 18 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1806946
string GDS_FILE /home/matt/work/asic-workshop/shuttle8/project5-walkthrough-mpw8/openlane/rgb_mixer/runs/23_01_03_13_12/results/signoff/rgb_mixer.magic.gds
string GDS_START 277910
<< end >>

