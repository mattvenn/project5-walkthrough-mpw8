// This is the unpowered netlist.
module rgb_mixer (clk,
    enc0_a,
    enc0_b,
    enc1_a,
    enc1_b,
    enc2_a,
    enc2_b,
    pwm0_out,
    pwm1_out,
    pwm2_out,
    reset,
    sync,
    io_oeb);
 input clk;
 input enc0_a;
 input enc0_b;
 input enc1_a;
 input enc1_b;
 input enc2_a;
 input enc2_b;
 output pwm0_out;
 output pwm1_out;
 output pwm2_out;
 input reset;
 output sync;
 output [3:0] io_oeb;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire _400_;
 wire _401_;
 wire _402_;
 wire _403_;
 wire _404_;
 wire _405_;
 wire _406_;
 wire _407_;
 wire _408_;
 wire _409_;
 wire _410_;
 wire _411_;
 wire _412_;
 wire _413_;
 wire _414_;
 wire _415_;
 wire _416_;
 wire _417_;
 wire _418_;
 wire _419_;
 wire _420_;
 wire _421_;
 wire _422_;
 wire _423_;
 wire _424_;
 wire _425_;
 wire \debounce0_a.button_hist[0] ;
 wire \debounce0_a.button_hist[1] ;
 wire \debounce0_a.button_hist[2] ;
 wire \debounce0_a.button_hist[3] ;
 wire \debounce0_a.button_hist[4] ;
 wire \debounce0_a.button_hist[5] ;
 wire \debounce0_a.button_hist[6] ;
 wire \debounce0_a.button_hist[7] ;
 wire \debounce0_a.debounced ;
 wire \debounce0_b.button_hist[0] ;
 wire \debounce0_b.button_hist[1] ;
 wire \debounce0_b.button_hist[2] ;
 wire \debounce0_b.button_hist[3] ;
 wire \debounce0_b.button_hist[4] ;
 wire \debounce0_b.button_hist[5] ;
 wire \debounce0_b.button_hist[6] ;
 wire \debounce0_b.button_hist[7] ;
 wire \debounce0_b.debounced ;
 wire \debounce1_a.button_hist[0] ;
 wire \debounce1_a.button_hist[1] ;
 wire \debounce1_a.button_hist[2] ;
 wire \debounce1_a.button_hist[3] ;
 wire \debounce1_a.button_hist[4] ;
 wire \debounce1_a.button_hist[5] ;
 wire \debounce1_a.button_hist[6] ;
 wire \debounce1_a.button_hist[7] ;
 wire \debounce1_a.debounced ;
 wire \debounce1_b.button_hist[0] ;
 wire \debounce1_b.button_hist[1] ;
 wire \debounce1_b.button_hist[2] ;
 wire \debounce1_b.button_hist[3] ;
 wire \debounce1_b.button_hist[4] ;
 wire \debounce1_b.button_hist[5] ;
 wire \debounce1_b.button_hist[6] ;
 wire \debounce1_b.button_hist[7] ;
 wire \debounce1_b.debounced ;
 wire \debounce2_a.button_hist[0] ;
 wire \debounce2_a.button_hist[1] ;
 wire \debounce2_a.button_hist[2] ;
 wire \debounce2_a.button_hist[3] ;
 wire \debounce2_a.button_hist[4] ;
 wire \debounce2_a.button_hist[5] ;
 wire \debounce2_a.button_hist[6] ;
 wire \debounce2_a.button_hist[7] ;
 wire \debounce2_a.debounced ;
 wire \debounce2_b.button_hist[0] ;
 wire \debounce2_b.button_hist[1] ;
 wire \debounce2_b.button_hist[2] ;
 wire \debounce2_b.button_hist[3] ;
 wire \debounce2_b.button_hist[4] ;
 wire \debounce2_b.button_hist[5] ;
 wire \debounce2_b.button_hist[6] ;
 wire \debounce2_b.button_hist[7] ;
 wire \debounce2_b.debounced ;
 wire \encoder0.old_a ;
 wire \encoder0.old_b ;
 wire \encoder0.value[0] ;
 wire \encoder0.value[1] ;
 wire \encoder0.value[2] ;
 wire \encoder0.value[3] ;
 wire \encoder0.value[4] ;
 wire \encoder0.value[5] ;
 wire \encoder0.value[6] ;
 wire \encoder0.value[7] ;
 wire \encoder1.old_a ;
 wire \encoder1.old_b ;
 wire \encoder1.value[0] ;
 wire \encoder1.value[1] ;
 wire \encoder1.value[2] ;
 wire \encoder1.value[3] ;
 wire \encoder1.value[4] ;
 wire \encoder1.value[5] ;
 wire \encoder1.value[6] ;
 wire \encoder1.value[7] ;
 wire \encoder2.old_a ;
 wire \encoder2.old_b ;
 wire \encoder2.value[0] ;
 wire \encoder2.value[1] ;
 wire \encoder2.value[2] ;
 wire \encoder2.value[3] ;
 wire \encoder2.value[4] ;
 wire \encoder2.value[5] ;
 wire \encoder2.value[6] ;
 wire \encoder2.value[7] ;
 wire net13;
 wire net14;
 wire net15;
 wire clknet_0_clk;
 wire \pwm0.count[0] ;
 wire \pwm0.count[1] ;
 wire \pwm0.count[2] ;
 wire \pwm0.count[3] ;
 wire \pwm0.count[4] ;
 wire \pwm0.count[5] ;
 wire \pwm0.count[6] ;
 wire \pwm0.count[7] ;
 wire \pwm1.count[0] ;
 wire \pwm1.count[1] ;
 wire \pwm1.count[2] ;
 wire \pwm1.count[3] ;
 wire \pwm1.count[4] ;
 wire \pwm1.count[5] ;
 wire \pwm1.count[6] ;
 wire \pwm1.count[7] ;
 wire \pwm2.count[0] ;
 wire \pwm2.count[1] ;
 wire \pwm2.count[2] ;
 wire \pwm2.count[3] ;
 wire \pwm2.count[4] ;
 wire \pwm2.count[5] ;
 wire \pwm2.count[6] ;
 wire \pwm2.count[7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;

 sky130_fd_sc_hd__clkinv_2 _426_ (.A(net7),
    .Y(_108_));
 sky130_fd_sc_hd__buf_2 _427_ (.A(_108_),
    .X(_109_));
 sky130_fd_sc_hd__or2b_1 _428_ (.A(\encoder0.value[7] ),
    .B_N(\pwm0.count[7] ),
    .X(_110_));
 sky130_fd_sc_hd__inv_2 _429_ (.A(\pwm0.count[7] ),
    .Y(_111_));
 sky130_fd_sc_hd__inv_2 _430_ (.A(\pwm0.count[6] ),
    .Y(_112_));
 sky130_fd_sc_hd__inv_2 _431_ (.A(\pwm0.count[5] ),
    .Y(_113_));
 sky130_fd_sc_hd__inv_2 _432_ (.A(\pwm0.count[4] ),
    .Y(_114_));
 sky130_fd_sc_hd__inv_2 _433_ (.A(\pwm0.count[3] ),
    .Y(_115_));
 sky130_fd_sc_hd__inv_2 _434_ (.A(\pwm0.count[2] ),
    .Y(_116_));
 sky130_fd_sc_hd__inv_2 _435_ (.A(\pwm0.count[1] ),
    .Y(_117_));
 sky130_fd_sc_hd__o22a_1 _436_ (.A1(\encoder0.value[2] ),
    .A2(_116_),
    .B1(_117_),
    .B2(\encoder0.value[1] ),
    .X(_118_));
 sky130_fd_sc_hd__inv_2 _437_ (.A(\pwm0.count[0] ),
    .Y(_119_));
 sky130_fd_sc_hd__o21ba_1 _438_ (.A1(\encoder0.value[0] ),
    .A2(_119_),
    .B1_N(_110_),
    .X(_120_));
 sky130_fd_sc_hd__a221o_1 _439_ (.A1(\encoder0.value[1] ),
    .A2(_117_),
    .B1(_119_),
    .B2(\encoder0.value[0] ),
    .C1(_120_),
    .X(_121_));
 sky130_fd_sc_hd__a22o_1 _440_ (.A1(\encoder0.value[3] ),
    .A2(_115_),
    .B1(_116_),
    .B2(\encoder0.value[2] ),
    .X(_122_));
 sky130_fd_sc_hd__a21o_1 _441_ (.A1(_118_),
    .A2(_121_),
    .B1(_122_),
    .X(_123_));
 sky130_fd_sc_hd__o221a_1 _442_ (.A1(\encoder0.value[4] ),
    .A2(_114_),
    .B1(_115_),
    .B2(\encoder0.value[3] ),
    .C1(_123_),
    .X(_124_));
 sky130_fd_sc_hd__a221o_1 _443_ (.A1(\encoder0.value[5] ),
    .A2(_113_),
    .B1(_114_),
    .B2(\encoder0.value[4] ),
    .C1(_124_),
    .X(_125_));
 sky130_fd_sc_hd__o221a_1 _444_ (.A1(\encoder0.value[6] ),
    .A2(_112_),
    .B1(_113_),
    .B2(\encoder0.value[5] ),
    .C1(_125_),
    .X(_126_));
 sky130_fd_sc_hd__a221o_1 _445_ (.A1(\encoder0.value[7] ),
    .A2(_111_),
    .B1(_112_),
    .B2(\encoder0.value[6] ),
    .C1(_126_),
    .X(_127_));
 sky130_fd_sc_hd__and3_1 _446_ (.A(_109_),
    .B(_110_),
    .C(_127_),
    .X(_128_));
 sky130_fd_sc_hd__clkbuf_1 _447_ (.A(_128_),
    .X(net8));
 sky130_fd_sc_hd__inv_2 _448_ (.A(\encoder1.value[7] ),
    .Y(_129_));
 sky130_fd_sc_hd__inv_2 _449_ (.A(\encoder1.value[6] ),
    .Y(_130_));
 sky130_fd_sc_hd__inv_2 _450_ (.A(\encoder1.value[5] ),
    .Y(_131_));
 sky130_fd_sc_hd__inv_2 _451_ (.A(\encoder1.value[4] ),
    .Y(_132_));
 sky130_fd_sc_hd__inv_2 _452_ (.A(\encoder1.value[3] ),
    .Y(_133_));
 sky130_fd_sc_hd__or2_1 _453_ (.A(_133_),
    .B(\pwm1.count[3] ),
    .X(_134_));
 sky130_fd_sc_hd__inv_2 _454_ (.A(\encoder1.value[2] ),
    .Y(_135_));
 sky130_fd_sc_hd__inv_2 _455_ (.A(\encoder1.value[1] ),
    .Y(_136_));
 sky130_fd_sc_hd__inv_2 _456_ (.A(\encoder1.value[0] ),
    .Y(_137_));
 sky130_fd_sc_hd__a211o_1 _457_ (.A1(_136_),
    .A2(\pwm1.count[1] ),
    .B1(\pwm1.count[0] ),
    .C1(_137_),
    .X(_138_));
 sky130_fd_sc_hd__o221a_1 _458_ (.A1(_135_),
    .A2(\pwm1.count[2] ),
    .B1(\pwm1.count[1] ),
    .B2(_136_),
    .C1(_138_),
    .X(_139_));
 sky130_fd_sc_hd__a221o_1 _459_ (.A1(_133_),
    .A2(\pwm1.count[3] ),
    .B1(\pwm1.count[2] ),
    .B2(_135_),
    .C1(_139_),
    .X(_140_));
 sky130_fd_sc_hd__a22o_1 _460_ (.A1(_132_),
    .A2(\pwm1.count[4] ),
    .B1(_134_),
    .B2(_140_),
    .X(_141_));
 sky130_fd_sc_hd__o221a_1 _461_ (.A1(_131_),
    .A2(\pwm1.count[5] ),
    .B1(\pwm1.count[4] ),
    .B2(_132_),
    .C1(_141_),
    .X(_142_));
 sky130_fd_sc_hd__a221o_1 _462_ (.A1(_130_),
    .A2(\pwm1.count[6] ),
    .B1(\pwm1.count[5] ),
    .B2(_131_),
    .C1(_142_),
    .X(_143_));
 sky130_fd_sc_hd__o221a_1 _463_ (.A1(_129_),
    .A2(\pwm1.count[7] ),
    .B1(\pwm1.count[6] ),
    .B2(_130_),
    .C1(_143_),
    .X(_144_));
 sky130_fd_sc_hd__clkbuf_4 _464_ (.A(net7),
    .X(_145_));
 sky130_fd_sc_hd__a211oi_1 _465_ (.A1(_129_),
    .A2(\pwm1.count[7] ),
    .B1(_144_),
    .C1(_145_),
    .Y(net9));
 sky130_fd_sc_hd__inv_2 _466_ (.A(\encoder2.value[7] ),
    .Y(_146_));
 sky130_fd_sc_hd__inv_2 _467_ (.A(\encoder2.value[6] ),
    .Y(_147_));
 sky130_fd_sc_hd__inv_2 _468_ (.A(\encoder2.value[5] ),
    .Y(_148_));
 sky130_fd_sc_hd__inv_2 _469_ (.A(\encoder2.value[4] ),
    .Y(_149_));
 sky130_fd_sc_hd__inv_2 _470_ (.A(\encoder2.value[3] ),
    .Y(_150_));
 sky130_fd_sc_hd__or2_1 _471_ (.A(_150_),
    .B(\pwm2.count[3] ),
    .X(_151_));
 sky130_fd_sc_hd__inv_2 _472_ (.A(\encoder2.value[2] ),
    .Y(_152_));
 sky130_fd_sc_hd__inv_2 _473_ (.A(\encoder2.value[1] ),
    .Y(_153_));
 sky130_fd_sc_hd__inv_2 _474_ (.A(\encoder2.value[0] ),
    .Y(_154_));
 sky130_fd_sc_hd__a211o_1 _475_ (.A1(_153_),
    .A2(\pwm2.count[1] ),
    .B1(\pwm2.count[0] ),
    .C1(_154_),
    .X(_155_));
 sky130_fd_sc_hd__o221a_1 _476_ (.A1(_152_),
    .A2(\pwm2.count[2] ),
    .B1(\pwm2.count[1] ),
    .B2(_153_),
    .C1(_155_),
    .X(_156_));
 sky130_fd_sc_hd__a221o_1 _477_ (.A1(_150_),
    .A2(\pwm2.count[3] ),
    .B1(\pwm2.count[2] ),
    .B2(_152_),
    .C1(_156_),
    .X(_157_));
 sky130_fd_sc_hd__a22o_1 _478_ (.A1(_149_),
    .A2(\pwm2.count[4] ),
    .B1(_151_),
    .B2(_157_),
    .X(_158_));
 sky130_fd_sc_hd__o221a_1 _479_ (.A1(_148_),
    .A2(\pwm2.count[5] ),
    .B1(\pwm2.count[4] ),
    .B2(_149_),
    .C1(_158_),
    .X(_159_));
 sky130_fd_sc_hd__a221o_1 _480_ (.A1(_147_),
    .A2(\pwm2.count[6] ),
    .B1(\pwm2.count[5] ),
    .B2(_148_),
    .C1(_159_),
    .X(_160_));
 sky130_fd_sc_hd__o221a_1 _481_ (.A1(_146_),
    .A2(\pwm2.count[7] ),
    .B1(\pwm2.count[6] ),
    .B2(_147_),
    .C1(_160_),
    .X(_161_));
 sky130_fd_sc_hd__a211oi_2 _482_ (.A1(_146_),
    .A2(\pwm2.count[7] ),
    .B1(_161_),
    .C1(_145_),
    .Y(net10));
 sky130_fd_sc_hd__clkbuf_4 _483_ (.A(_109_),
    .X(_162_));
 sky130_fd_sc_hd__and4_1 _484_ (.A(\debounce0_a.button_hist[5] ),
    .B(\debounce0_a.button_hist[4] ),
    .C(\debounce0_a.button_hist[7] ),
    .D(\debounce0_a.button_hist[6] ),
    .X(_163_));
 sky130_fd_sc_hd__and4_1 _485_ (.A(\debounce0_a.button_hist[1] ),
    .B(\debounce0_a.button_hist[0] ),
    .C(\debounce0_a.button_hist[3] ),
    .D(\debounce0_a.button_hist[2] ),
    .X(_164_));
 sky130_fd_sc_hd__or4_1 _486_ (.A(\debounce0_a.button_hist[1] ),
    .B(\debounce0_a.button_hist[0] ),
    .C(\debounce0_a.button_hist[3] ),
    .D(\debounce0_a.button_hist[2] ),
    .X(_165_));
 sky130_fd_sc_hd__or4_1 _487_ (.A(\debounce0_a.button_hist[5] ),
    .B(\debounce0_a.button_hist[4] ),
    .C(\debounce0_a.button_hist[7] ),
    .D(\debounce0_a.button_hist[6] ),
    .X(_166_));
 sky130_fd_sc_hd__or2_1 _488_ (.A(_165_),
    .B(_166_),
    .X(_167_));
 sky130_fd_sc_hd__and2_1 _489_ (.A(\debounce0_a.debounced ),
    .B(_108_),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_1 _490_ (.A(_168_),
    .X(_054_));
 sky130_fd_sc_hd__a32o_1 _491_ (.A1(_162_),
    .A2(_163_),
    .A3(_164_),
    .B1(_167_),
    .B2(_054_),
    .X(_000_));
 sky130_fd_sc_hd__clkbuf_4 _492_ (.A(_108_),
    .X(_169_));
 sky130_fd_sc_hd__and2_1 _493_ (.A(_169_),
    .B(net1),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_1 _494_ (.A(_170_),
    .X(_001_));
 sky130_fd_sc_hd__and2_1 _495_ (.A(\debounce0_a.button_hist[0] ),
    .B(_169_),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _496_ (.A(_171_),
    .X(_002_));
 sky130_fd_sc_hd__clkbuf_2 _497_ (.A(_109_),
    .X(_172_));
 sky130_fd_sc_hd__and2_1 _498_ (.A(\debounce0_a.button_hist[1] ),
    .B(_172_),
    .X(_173_));
 sky130_fd_sc_hd__clkbuf_1 _499_ (.A(_173_),
    .X(_003_));
 sky130_fd_sc_hd__and2_1 _500_ (.A(\debounce0_a.button_hist[2] ),
    .B(_169_),
    .X(_174_));
 sky130_fd_sc_hd__clkbuf_1 _501_ (.A(_174_),
    .X(_004_));
 sky130_fd_sc_hd__and2_1 _502_ (.A(\debounce0_a.button_hist[3] ),
    .B(_172_),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _503_ (.A(_175_),
    .X(_005_));
 sky130_fd_sc_hd__and2_1 _504_ (.A(\debounce0_a.button_hist[4] ),
    .B(_172_),
    .X(_176_));
 sky130_fd_sc_hd__clkbuf_1 _505_ (.A(_176_),
    .X(_006_));
 sky130_fd_sc_hd__and2_1 _506_ (.A(\debounce0_a.button_hist[5] ),
    .B(_172_),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _507_ (.A(_177_),
    .X(_007_));
 sky130_fd_sc_hd__and2_1 _508_ (.A(\debounce0_a.button_hist[6] ),
    .B(_172_),
    .X(_178_));
 sky130_fd_sc_hd__clkbuf_1 _509_ (.A(_178_),
    .X(_008_));
 sky130_fd_sc_hd__and2_1 _510_ (.A(\debounce0_b.button_hist[0] ),
    .B(_108_),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _511_ (.A(_179_),
    .X(_011_));
 sky130_fd_sc_hd__and4_1 _512_ (.A(\debounce0_b.button_hist[5] ),
    .B(\debounce0_b.button_hist[4] ),
    .C(\debounce0_b.button_hist[7] ),
    .D(\debounce0_b.button_hist[6] ),
    .X(_180_));
 sky130_fd_sc_hd__and3_1 _513_ (.A(\debounce0_b.button_hist[1] ),
    .B(\debounce0_b.button_hist[2] ),
    .C(_180_),
    .X(_181_));
 sky130_fd_sc_hd__or3_1 _514_ (.A(\debounce0_b.button_hist[1] ),
    .B(\debounce0_b.button_hist[0] ),
    .C(\debounce0_b.button_hist[3] ),
    .X(_182_));
 sky130_fd_sc_hd__or4_1 _515_ (.A(\debounce0_b.button_hist[5] ),
    .B(\debounce0_b.button_hist[4] ),
    .C(\debounce0_b.button_hist[7] ),
    .D(\debounce0_b.button_hist[6] ),
    .X(_183_));
 sky130_fd_sc_hd__o31a_1 _516_ (.A1(\debounce0_b.button_hist[2] ),
    .A2(_182_),
    .A3(_183_),
    .B1(\debounce0_b.debounced ),
    .X(_184_));
 sky130_fd_sc_hd__a32o_1 _517_ (.A1(\debounce0_b.button_hist[3] ),
    .A2(_011_),
    .A3(_181_),
    .B1(_162_),
    .B2(_184_),
    .X(_009_));
 sky130_fd_sc_hd__and2_1 _518_ (.A(_169_),
    .B(net2),
    .X(_185_));
 sky130_fd_sc_hd__clkbuf_1 _519_ (.A(_185_),
    .X(_010_));
 sky130_fd_sc_hd__and2_1 _520_ (.A(\debounce0_b.button_hist[1] ),
    .B(_172_),
    .X(_186_));
 sky130_fd_sc_hd__clkbuf_1 _521_ (.A(_186_),
    .X(_012_));
 sky130_fd_sc_hd__and2_1 _522_ (.A(\debounce0_b.button_hist[2] ),
    .B(_172_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_1 _523_ (.A(_187_),
    .X(_013_));
 sky130_fd_sc_hd__and2_1 _524_ (.A(\debounce0_b.button_hist[3] ),
    .B(_172_),
    .X(_188_));
 sky130_fd_sc_hd__clkbuf_1 _525_ (.A(_188_),
    .X(_014_));
 sky130_fd_sc_hd__and2_1 _526_ (.A(\debounce0_b.button_hist[4] ),
    .B(_172_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _527_ (.A(_189_),
    .X(_015_));
 sky130_fd_sc_hd__clkbuf_2 _528_ (.A(_109_),
    .X(_190_));
 sky130_fd_sc_hd__and2_1 _529_ (.A(\debounce0_b.button_hist[5] ),
    .B(_190_),
    .X(_191_));
 sky130_fd_sc_hd__clkbuf_1 _530_ (.A(_191_),
    .X(_016_));
 sky130_fd_sc_hd__and2_1 _531_ (.A(\debounce0_b.button_hist[6] ),
    .B(_190_),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _532_ (.A(_192_),
    .X(_017_));
 sky130_fd_sc_hd__and2_1 _533_ (.A(\debounce1_a.button_hist[0] ),
    .B(_108_),
    .X(_193_));
 sky130_fd_sc_hd__clkbuf_1 _534_ (.A(_193_),
    .X(_020_));
 sky130_fd_sc_hd__and4_1 _535_ (.A(\debounce1_a.button_hist[5] ),
    .B(\debounce1_a.button_hist[4] ),
    .C(\debounce1_a.button_hist[7] ),
    .D(\debounce1_a.button_hist[6] ),
    .X(_194_));
 sky130_fd_sc_hd__and3_1 _536_ (.A(\debounce1_a.button_hist[1] ),
    .B(\debounce1_a.button_hist[2] ),
    .C(_194_),
    .X(_195_));
 sky130_fd_sc_hd__or3_1 _537_ (.A(\debounce1_a.button_hist[1] ),
    .B(\debounce1_a.button_hist[0] ),
    .C(\debounce1_a.button_hist[3] ),
    .X(_196_));
 sky130_fd_sc_hd__or4_1 _538_ (.A(\debounce1_a.button_hist[5] ),
    .B(\debounce1_a.button_hist[4] ),
    .C(\debounce1_a.button_hist[7] ),
    .D(\debounce1_a.button_hist[6] ),
    .X(_197_));
 sky130_fd_sc_hd__o31a_1 _539_ (.A1(\debounce1_a.button_hist[2] ),
    .A2(_196_),
    .A3(_197_),
    .B1(\debounce1_a.debounced ),
    .X(_198_));
 sky130_fd_sc_hd__a32o_1 _540_ (.A1(\debounce1_a.button_hist[3] ),
    .A2(_020_),
    .A3(_195_),
    .B1(_162_),
    .B2(_198_),
    .X(_018_));
 sky130_fd_sc_hd__and2_1 _541_ (.A(_169_),
    .B(net3),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _542_ (.A(_199_),
    .X(_019_));
 sky130_fd_sc_hd__and2_1 _543_ (.A(\debounce1_a.button_hist[1] ),
    .B(_190_),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _544_ (.A(_200_),
    .X(_021_));
 sky130_fd_sc_hd__and2_1 _545_ (.A(\debounce1_a.button_hist[2] ),
    .B(_190_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _546_ (.A(_201_),
    .X(_022_));
 sky130_fd_sc_hd__and2_1 _547_ (.A(\debounce1_a.button_hist[3] ),
    .B(_190_),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _548_ (.A(_202_),
    .X(_023_));
 sky130_fd_sc_hd__and2_1 _549_ (.A(\debounce1_a.button_hist[4] ),
    .B(_190_),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _550_ (.A(_203_),
    .X(_024_));
 sky130_fd_sc_hd__and2_1 _551_ (.A(\debounce1_a.button_hist[5] ),
    .B(_190_),
    .X(_204_));
 sky130_fd_sc_hd__clkbuf_1 _552_ (.A(_204_),
    .X(_025_));
 sky130_fd_sc_hd__and2_1 _553_ (.A(\debounce1_a.button_hist[6] ),
    .B(_190_),
    .X(_205_));
 sky130_fd_sc_hd__clkbuf_1 _554_ (.A(_205_),
    .X(_026_));
 sky130_fd_sc_hd__and2_1 _555_ (.A(\debounce1_b.button_hist[0] ),
    .B(_108_),
    .X(_206_));
 sky130_fd_sc_hd__clkbuf_1 _556_ (.A(_206_),
    .X(_029_));
 sky130_fd_sc_hd__and4_1 _557_ (.A(\debounce1_b.button_hist[5] ),
    .B(\debounce1_b.button_hist[4] ),
    .C(\debounce1_b.button_hist[7] ),
    .D(\debounce1_b.button_hist[6] ),
    .X(_207_));
 sky130_fd_sc_hd__and3_1 _558_ (.A(\debounce1_b.button_hist[1] ),
    .B(\debounce1_b.button_hist[2] ),
    .C(_207_),
    .X(_208_));
 sky130_fd_sc_hd__or4_1 _559_ (.A(\debounce1_b.button_hist[1] ),
    .B(\debounce1_b.button_hist[0] ),
    .C(\debounce1_b.button_hist[3] ),
    .D(\debounce1_b.button_hist[2] ),
    .X(_209_));
 sky130_fd_sc_hd__or4_1 _560_ (.A(\debounce1_b.button_hist[5] ),
    .B(\debounce1_b.button_hist[4] ),
    .C(\debounce1_b.button_hist[7] ),
    .D(\debounce1_b.button_hist[6] ),
    .X(_210_));
 sky130_fd_sc_hd__o211a_1 _561_ (.A1(_209_),
    .A2(_210_),
    .B1(\debounce1_b.debounced ),
    .C1(_109_),
    .X(_211_));
 sky130_fd_sc_hd__a31o_1 _562_ (.A1(\debounce1_b.button_hist[3] ),
    .A2(_029_),
    .A3(_208_),
    .B1(_211_),
    .X(_027_));
 sky130_fd_sc_hd__and2_1 _563_ (.A(_169_),
    .B(net4),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _564_ (.A(_212_),
    .X(_028_));
 sky130_fd_sc_hd__clkbuf_2 _565_ (.A(_109_),
    .X(_213_));
 sky130_fd_sc_hd__and2_1 _566_ (.A(\debounce1_b.button_hist[1] ),
    .B(_213_),
    .X(_214_));
 sky130_fd_sc_hd__clkbuf_1 _567_ (.A(_214_),
    .X(_030_));
 sky130_fd_sc_hd__and2_1 _568_ (.A(\debounce1_b.button_hist[2] ),
    .B(_213_),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _569_ (.A(_215_),
    .X(_031_));
 sky130_fd_sc_hd__and2_1 _570_ (.A(\debounce1_b.button_hist[3] ),
    .B(_213_),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _571_ (.A(_216_),
    .X(_032_));
 sky130_fd_sc_hd__and2_1 _572_ (.A(\debounce1_b.button_hist[4] ),
    .B(_213_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _573_ (.A(_217_),
    .X(_033_));
 sky130_fd_sc_hd__and2_1 _574_ (.A(\debounce1_b.button_hist[5] ),
    .B(_213_),
    .X(_218_));
 sky130_fd_sc_hd__clkbuf_1 _575_ (.A(_218_),
    .X(_034_));
 sky130_fd_sc_hd__and2_1 _576_ (.A(\debounce1_b.button_hist[6] ),
    .B(_213_),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_1 _577_ (.A(_219_),
    .X(_035_));
 sky130_fd_sc_hd__clkbuf_4 _578_ (.A(_109_),
    .X(_220_));
 sky130_fd_sc_hd__and4_1 _579_ (.A(\debounce2_a.button_hist[5] ),
    .B(\debounce2_a.button_hist[4] ),
    .C(\debounce2_a.button_hist[7] ),
    .D(\debounce2_a.button_hist[6] ),
    .X(_221_));
 sky130_fd_sc_hd__and4_1 _580_ (.A(\debounce2_a.button_hist[1] ),
    .B(\debounce2_a.button_hist[0] ),
    .C(\debounce2_a.button_hist[3] ),
    .D(\debounce2_a.button_hist[2] ),
    .X(_222_));
 sky130_fd_sc_hd__or4_1 _581_ (.A(\debounce2_a.button_hist[5] ),
    .B(\debounce2_a.button_hist[4] ),
    .C(\debounce2_a.button_hist[7] ),
    .D(\debounce2_a.button_hist[6] ),
    .X(_223_));
 sky130_fd_sc_hd__or3_1 _582_ (.A(\debounce2_a.button_hist[3] ),
    .B(\debounce2_a.button_hist[2] ),
    .C(_223_),
    .X(_224_));
 sky130_fd_sc_hd__and2_1 _583_ (.A(\debounce2_a.debounced ),
    .B(_108_),
    .X(_225_));
 sky130_fd_sc_hd__clkbuf_1 _584_ (.A(_225_),
    .X(_081_));
 sky130_fd_sc_hd__o31a_1 _585_ (.A1(\debounce2_a.button_hist[1] ),
    .A2(\debounce2_a.button_hist[0] ),
    .A3(_224_),
    .B1(_081_),
    .X(_226_));
 sky130_fd_sc_hd__a31o_1 _586_ (.A1(_220_),
    .A2(_221_),
    .A3(_222_),
    .B1(_226_),
    .X(_036_));
 sky130_fd_sc_hd__and2_1 _587_ (.A(_169_),
    .B(net5),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _588_ (.A(_227_),
    .X(_037_));
 sky130_fd_sc_hd__and2_1 _589_ (.A(\debounce2_a.button_hist[0] ),
    .B(_213_),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_1 _590_ (.A(_228_),
    .X(_038_));
 sky130_fd_sc_hd__and2_1 _591_ (.A(\debounce2_a.button_hist[1] ),
    .B(_213_),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _592_ (.A(_229_),
    .X(_039_));
 sky130_fd_sc_hd__and2_1 _593_ (.A(\debounce2_a.button_hist[2] ),
    .B(_213_),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _594_ (.A(_230_),
    .X(_040_));
 sky130_fd_sc_hd__and2_1 _595_ (.A(\debounce2_a.button_hist[3] ),
    .B(_213_),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_1 _596_ (.A(_231_),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_2 _597_ (.A(_109_),
    .X(_232_));
 sky130_fd_sc_hd__and2_1 _598_ (.A(\debounce2_a.button_hist[4] ),
    .B(_232_),
    .X(_233_));
 sky130_fd_sc_hd__clkbuf_1 _599_ (.A(_233_),
    .X(_042_));
 sky130_fd_sc_hd__and2_1 _600_ (.A(\debounce2_a.button_hist[5] ),
    .B(_232_),
    .X(_234_));
 sky130_fd_sc_hd__clkbuf_1 _601_ (.A(_234_),
    .X(_043_));
 sky130_fd_sc_hd__and2_1 _602_ (.A(\debounce2_a.button_hist[6] ),
    .B(_232_),
    .X(_235_));
 sky130_fd_sc_hd__clkbuf_1 _603_ (.A(_235_),
    .X(_044_));
 sky130_fd_sc_hd__and2_1 _604_ (.A(\debounce2_b.button_hist[1] ),
    .B(_108_),
    .X(_236_));
 sky130_fd_sc_hd__clkbuf_1 _605_ (.A(_236_),
    .X(_057_));
 sky130_fd_sc_hd__and4_1 _606_ (.A(\debounce2_b.button_hist[5] ),
    .B(\debounce2_b.button_hist[4] ),
    .C(\debounce2_b.button_hist[7] ),
    .D(\debounce2_b.button_hist[6] ),
    .X(_237_));
 sky130_fd_sc_hd__and3_1 _607_ (.A(\debounce2_b.button_hist[0] ),
    .B(\debounce2_b.button_hist[3] ),
    .C(_237_),
    .X(_238_));
 sky130_fd_sc_hd__or4_1 _608_ (.A(\debounce2_b.button_hist[1] ),
    .B(\debounce2_b.button_hist[0] ),
    .C(\debounce2_b.button_hist[3] ),
    .D(\debounce2_b.button_hist[2] ),
    .X(_239_));
 sky130_fd_sc_hd__or4_1 _609_ (.A(\debounce2_b.button_hist[5] ),
    .B(\debounce2_b.button_hist[4] ),
    .C(\debounce2_b.button_hist[7] ),
    .D(\debounce2_b.button_hist[6] ),
    .X(_240_));
 sky130_fd_sc_hd__o211a_1 _610_ (.A1(_239_),
    .A2(_240_),
    .B1(\debounce2_b.debounced ),
    .C1(_109_),
    .X(_241_));
 sky130_fd_sc_hd__a31o_1 _611_ (.A1(\debounce2_b.button_hist[2] ),
    .A2(_057_),
    .A3(_238_),
    .B1(_241_),
    .X(_045_));
 sky130_fd_sc_hd__nor2_1 _612_ (.A(_145_),
    .B(\pwm2.count[0] ),
    .Y(_046_));
 sky130_fd_sc_hd__clkbuf_4 _613_ (.A(net7),
    .X(_242_));
 sky130_fd_sc_hd__a21oi_1 _614_ (.A1(\pwm2.count[1] ),
    .A2(\pwm2.count[0] ),
    .B1(_242_),
    .Y(_243_));
 sky130_fd_sc_hd__o21a_1 _615_ (.A1(\pwm2.count[1] ),
    .A2(\pwm2.count[0] ),
    .B1(_243_),
    .X(_047_));
 sky130_fd_sc_hd__a21oi_1 _616_ (.A1(\pwm2.count[1] ),
    .A2(\pwm2.count[0] ),
    .B1(\pwm2.count[2] ),
    .Y(_244_));
 sky130_fd_sc_hd__and3_1 _617_ (.A(\pwm2.count[2] ),
    .B(\pwm2.count[1] ),
    .C(\pwm2.count[0] ),
    .X(_245_));
 sky130_fd_sc_hd__nor3_1 _618_ (.A(_145_),
    .B(_244_),
    .C(_245_),
    .Y(_048_));
 sky130_fd_sc_hd__and2_1 _619_ (.A(\pwm2.count[3] ),
    .B(_245_),
    .X(_246_));
 sky130_fd_sc_hd__o21ai_1 _620_ (.A1(\pwm2.count[3] ),
    .A2(_245_),
    .B1(_162_),
    .Y(_247_));
 sky130_fd_sc_hd__nor2_1 _621_ (.A(_246_),
    .B(_247_),
    .Y(_049_));
 sky130_fd_sc_hd__and3_1 _622_ (.A(\pwm2.count[4] ),
    .B(\pwm2.count[3] ),
    .C(_245_),
    .X(_248_));
 sky130_fd_sc_hd__o21ai_1 _623_ (.A1(\pwm2.count[4] ),
    .A2(_246_),
    .B1(_162_),
    .Y(_249_));
 sky130_fd_sc_hd__nor2_1 _624_ (.A(_248_),
    .B(_249_),
    .Y(_050_));
 sky130_fd_sc_hd__and2_1 _625_ (.A(\pwm2.count[5] ),
    .B(_248_),
    .X(_250_));
 sky130_fd_sc_hd__nor2_1 _626_ (.A(_242_),
    .B(_250_),
    .Y(_251_));
 sky130_fd_sc_hd__o21a_1 _627_ (.A1(\pwm2.count[5] ),
    .A2(_248_),
    .B1(_251_),
    .X(_051_));
 sky130_fd_sc_hd__and3_1 _628_ (.A(\pwm2.count[6] ),
    .B(\pwm2.count[5] ),
    .C(_248_),
    .X(_252_));
 sky130_fd_sc_hd__o21ai_1 _629_ (.A1(\pwm2.count[6] ),
    .A2(_250_),
    .B1(_162_),
    .Y(_253_));
 sky130_fd_sc_hd__nor2_1 _630_ (.A(_252_),
    .B(_253_),
    .Y(_052_));
 sky130_fd_sc_hd__a21oi_1 _631_ (.A1(\pwm2.count[7] ),
    .A2(_252_),
    .B1(_242_),
    .Y(_254_));
 sky130_fd_sc_hd__o21a_1 _632_ (.A1(\pwm2.count[7] ),
    .A2(_252_),
    .B1(_254_),
    .X(_053_));
 sky130_fd_sc_hd__and2_1 _633_ (.A(_169_),
    .B(net6),
    .X(_255_));
 sky130_fd_sc_hd__clkbuf_1 _634_ (.A(_255_),
    .X(_055_));
 sky130_fd_sc_hd__and2_1 _635_ (.A(\debounce2_b.button_hist[0] ),
    .B(_232_),
    .X(_256_));
 sky130_fd_sc_hd__clkbuf_1 _636_ (.A(_256_),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _637_ (.A(\debounce2_b.button_hist[2] ),
    .B(_232_),
    .X(_257_));
 sky130_fd_sc_hd__clkbuf_1 _638_ (.A(_257_),
    .X(_058_));
 sky130_fd_sc_hd__and2_1 _639_ (.A(\debounce2_b.button_hist[3] ),
    .B(_232_),
    .X(_258_));
 sky130_fd_sc_hd__clkbuf_1 _640_ (.A(_258_),
    .X(_059_));
 sky130_fd_sc_hd__and2_1 _641_ (.A(\debounce2_b.button_hist[4] ),
    .B(_232_),
    .X(_259_));
 sky130_fd_sc_hd__clkbuf_1 _642_ (.A(_259_),
    .X(_060_));
 sky130_fd_sc_hd__and2_1 _643_ (.A(\debounce2_b.button_hist[5] ),
    .B(_232_),
    .X(_260_));
 sky130_fd_sc_hd__clkbuf_1 _644_ (.A(_260_),
    .X(_061_));
 sky130_fd_sc_hd__and2_1 _645_ (.A(\debounce2_b.button_hist[6] ),
    .B(_232_),
    .X(_261_));
 sky130_fd_sc_hd__clkbuf_1 _646_ (.A(_261_),
    .X(_062_));
 sky130_fd_sc_hd__and2b_1 _647_ (.A_N(\debounce0_a.debounced ),
    .B(\debounce0_b.debounced ),
    .X(_262_));
 sky130_fd_sc_hd__and2b_1 _648_ (.A_N(\debounce0_b.debounced ),
    .B(\debounce0_a.debounced ),
    .X(_263_));
 sky130_fd_sc_hd__and2_1 _649_ (.A(\encoder0.old_b ),
    .B(\encoder0.old_a ),
    .X(_264_));
 sky130_fd_sc_hd__nor2_1 _650_ (.A(\encoder0.old_b ),
    .B(\encoder0.old_a ),
    .Y(_265_));
 sky130_fd_sc_hd__o22a_2 _651_ (.A1(_262_),
    .A2(_263_),
    .B1(_264_),
    .B2(_265_),
    .X(_266_));
 sky130_fd_sc_hd__buf_2 _652_ (.A(_266_),
    .X(_267_));
 sky130_fd_sc_hd__a21oi_1 _653_ (.A1(\encoder0.value[0] ),
    .A2(_266_),
    .B1(_242_),
    .Y(_268_));
 sky130_fd_sc_hd__o21a_1 _654_ (.A1(\encoder0.value[0] ),
    .A2(_267_),
    .B1(_268_),
    .X(_063_));
 sky130_fd_sc_hd__o22a_1 _655_ (.A1(_262_),
    .A2(_264_),
    .B1(_265_),
    .B2(_263_),
    .X(_269_));
 sky130_fd_sc_hd__or2_1 _656_ (.A(\encoder0.value[1] ),
    .B(_269_),
    .X(_270_));
 sky130_fd_sc_hd__nand2_1 _657_ (.A(\encoder0.value[1] ),
    .B(_269_),
    .Y(_271_));
 sky130_fd_sc_hd__a21oi_1 _658_ (.A1(_270_),
    .A2(_271_),
    .B1(\encoder0.value[0] ),
    .Y(_272_));
 sky130_fd_sc_hd__and3_1 _659_ (.A(\encoder0.value[0] ),
    .B(_270_),
    .C(_271_),
    .X(_273_));
 sky130_fd_sc_hd__o21ai_1 _660_ (.A1(_272_),
    .A2(_273_),
    .B1(_266_),
    .Y(_274_));
 sky130_fd_sc_hd__clkbuf_4 _661_ (.A(_109_),
    .X(_275_));
 sky130_fd_sc_hd__o211a_1 _662_ (.A1(\encoder0.value[1] ),
    .A2(_267_),
    .B1(_274_),
    .C1(_275_),
    .X(_064_));
 sky130_fd_sc_hd__a21boi_1 _663_ (.A1(\encoder0.value[0] ),
    .A2(_270_),
    .B1_N(_271_),
    .Y(_276_));
 sky130_fd_sc_hd__or2_1 _664_ (.A(\encoder0.value[2] ),
    .B(_269_),
    .X(_277_));
 sky130_fd_sc_hd__clkbuf_4 _665_ (.A(_269_),
    .X(_278_));
 sky130_fd_sc_hd__nand2_1 _666_ (.A(\encoder0.value[2] ),
    .B(_278_),
    .Y(_279_));
 sky130_fd_sc_hd__nand2_1 _667_ (.A(_277_),
    .B(_279_),
    .Y(_280_));
 sky130_fd_sc_hd__xnor2_1 _668_ (.A(_276_),
    .B(_280_),
    .Y(_281_));
 sky130_fd_sc_hd__nand2_1 _669_ (.A(_267_),
    .B(_281_),
    .Y(_282_));
 sky130_fd_sc_hd__o211a_1 _670_ (.A1(\encoder0.value[2] ),
    .A2(_267_),
    .B1(_282_),
    .C1(_275_),
    .X(_065_));
 sky130_fd_sc_hd__xnor2_1 _671_ (.A(\encoder0.value[3] ),
    .B(_278_),
    .Y(_283_));
 sky130_fd_sc_hd__o21ai_1 _672_ (.A1(_276_),
    .A2(_280_),
    .B1(_279_),
    .Y(_284_));
 sky130_fd_sc_hd__a21boi_1 _673_ (.A1(_283_),
    .A2(_284_),
    .B1_N(_266_),
    .Y(_285_));
 sky130_fd_sc_hd__o21ai_1 _674_ (.A1(_283_),
    .A2(_284_),
    .B1(_285_),
    .Y(_286_));
 sky130_fd_sc_hd__o211a_1 _675_ (.A1(\encoder0.value[3] ),
    .A2(_267_),
    .B1(_286_),
    .C1(_275_),
    .X(_066_));
 sky130_fd_sc_hd__o21ai_1 _676_ (.A1(\encoder0.value[3] ),
    .A2(\encoder0.value[2] ),
    .B1(_278_),
    .Y(_287_));
 sky130_fd_sc_hd__o31a_1 _677_ (.A1(_276_),
    .A2(_280_),
    .A3(_283_),
    .B1(_287_),
    .X(_288_));
 sky130_fd_sc_hd__xnor2_1 _678_ (.A(\encoder0.value[4] ),
    .B(_278_),
    .Y(_289_));
 sky130_fd_sc_hd__and2_1 _679_ (.A(_288_),
    .B(_289_),
    .X(_290_));
 sky130_fd_sc_hd__nor2_1 _680_ (.A(_288_),
    .B(_289_),
    .Y(_291_));
 sky130_fd_sc_hd__o21ai_1 _681_ (.A1(_290_),
    .A2(_291_),
    .B1(_266_),
    .Y(_292_));
 sky130_fd_sc_hd__o211a_1 _682_ (.A1(\encoder0.value[4] ),
    .A2(_267_),
    .B1(_292_),
    .C1(_275_),
    .X(_067_));
 sky130_fd_sc_hd__xnor2_1 _683_ (.A(\encoder0.value[5] ),
    .B(_278_),
    .Y(_293_));
 sky130_fd_sc_hd__a21oi_1 _684_ (.A1(\encoder0.value[4] ),
    .A2(_278_),
    .B1(_291_),
    .Y(_294_));
 sky130_fd_sc_hd__xnor2_1 _685_ (.A(_293_),
    .B(_294_),
    .Y(_295_));
 sky130_fd_sc_hd__nor2_1 _686_ (.A(\encoder0.value[5] ),
    .B(_266_),
    .Y(_296_));
 sky130_fd_sc_hd__a211oi_1 _687_ (.A1(_267_),
    .A2(_295_),
    .B1(_296_),
    .C1(_145_),
    .Y(_068_));
 sky130_fd_sc_hd__nor2_1 _688_ (.A(\encoder0.value[6] ),
    .B(_278_),
    .Y(_297_));
 sky130_fd_sc_hd__nand2_1 _689_ (.A(\encoder0.value[6] ),
    .B(_278_),
    .Y(_298_));
 sky130_fd_sc_hd__or2b_1 _690_ (.A(_297_),
    .B_N(_298_),
    .X(_299_));
 sky130_fd_sc_hd__o21ai_1 _691_ (.A1(\encoder0.value[5] ),
    .A2(\encoder0.value[4] ),
    .B1(_278_),
    .Y(_300_));
 sky130_fd_sc_hd__o31a_1 _692_ (.A1(_288_),
    .A2(_289_),
    .A3(_293_),
    .B1(_300_),
    .X(_301_));
 sky130_fd_sc_hd__xnor2_1 _693_ (.A(_299_),
    .B(_301_),
    .Y(_302_));
 sky130_fd_sc_hd__nand2_1 _694_ (.A(_267_),
    .B(_302_),
    .Y(_303_));
 sky130_fd_sc_hd__o211a_1 _695_ (.A1(\encoder0.value[6] ),
    .A2(_267_),
    .B1(_303_),
    .C1(_275_),
    .X(_069_));
 sky130_fd_sc_hd__o21ai_1 _696_ (.A1(_297_),
    .A2(_301_),
    .B1(_298_),
    .Y(_304_));
 sky130_fd_sc_hd__xnor2_1 _697_ (.A(\encoder0.value[7] ),
    .B(_278_),
    .Y(_305_));
 sky130_fd_sc_hd__nor2_1 _698_ (.A(_304_),
    .B(_305_),
    .Y(_306_));
 sky130_fd_sc_hd__a21bo_1 _699_ (.A1(_304_),
    .A2(_305_),
    .B1_N(_266_),
    .X(_307_));
 sky130_fd_sc_hd__o221a_1 _700_ (.A1(\encoder0.value[7] ),
    .A2(_267_),
    .B1(_306_),
    .B2(_307_),
    .C1(_220_),
    .X(_070_));
 sky130_fd_sc_hd__and2_1 _701_ (.A(\debounce1_a.debounced ),
    .B(_190_),
    .X(_308_));
 sky130_fd_sc_hd__clkbuf_1 _702_ (.A(_308_),
    .X(_071_));
 sky130_fd_sc_hd__and2_1 _703_ (.A(\debounce0_b.debounced ),
    .B(_172_),
    .X(_309_));
 sky130_fd_sc_hd__clkbuf_1 _704_ (.A(_309_),
    .X(_072_));
 sky130_fd_sc_hd__and2b_1 _705_ (.A_N(\debounce1_a.debounced ),
    .B(\debounce1_b.debounced ),
    .X(_310_));
 sky130_fd_sc_hd__and2b_1 _706_ (.A_N(\debounce1_b.debounced ),
    .B(\debounce1_a.debounced ),
    .X(_311_));
 sky130_fd_sc_hd__and2_1 _707_ (.A(\encoder1.old_b ),
    .B(\encoder1.old_a ),
    .X(_312_));
 sky130_fd_sc_hd__nor2_1 _708_ (.A(\encoder1.old_b ),
    .B(\encoder1.old_a ),
    .Y(_313_));
 sky130_fd_sc_hd__o22a_2 _709_ (.A1(_310_),
    .A2(_311_),
    .B1(_312_),
    .B2(_313_),
    .X(_314_));
 sky130_fd_sc_hd__buf_2 _710_ (.A(_314_),
    .X(_315_));
 sky130_fd_sc_hd__a21oi_1 _711_ (.A1(\encoder1.value[0] ),
    .A2(_314_),
    .B1(_242_),
    .Y(_316_));
 sky130_fd_sc_hd__o21a_1 _712_ (.A1(\encoder1.value[0] ),
    .A2(_315_),
    .B1(_316_),
    .X(_073_));
 sky130_fd_sc_hd__o22a_1 _713_ (.A1(_310_),
    .A2(_312_),
    .B1(_313_),
    .B2(_311_),
    .X(_317_));
 sky130_fd_sc_hd__or2_1 _714_ (.A(\encoder1.value[1] ),
    .B(_317_),
    .X(_318_));
 sky130_fd_sc_hd__nand2_1 _715_ (.A(\encoder1.value[1] ),
    .B(_317_),
    .Y(_319_));
 sky130_fd_sc_hd__a21oi_1 _716_ (.A1(_318_),
    .A2(_319_),
    .B1(\encoder1.value[0] ),
    .Y(_320_));
 sky130_fd_sc_hd__and3_1 _717_ (.A(\encoder1.value[0] ),
    .B(_318_),
    .C(_319_),
    .X(_321_));
 sky130_fd_sc_hd__o21ai_1 _718_ (.A1(_320_),
    .A2(_321_),
    .B1(_314_),
    .Y(_322_));
 sky130_fd_sc_hd__o211a_1 _719_ (.A1(\encoder1.value[1] ),
    .A2(_315_),
    .B1(_322_),
    .C1(_275_),
    .X(_074_));
 sky130_fd_sc_hd__a21boi_1 _720_ (.A1(\encoder1.value[0] ),
    .A2(_318_),
    .B1_N(_319_),
    .Y(_323_));
 sky130_fd_sc_hd__or2_1 _721_ (.A(\encoder1.value[2] ),
    .B(_317_),
    .X(_324_));
 sky130_fd_sc_hd__clkbuf_4 _722_ (.A(_317_),
    .X(_325_));
 sky130_fd_sc_hd__nand2_1 _723_ (.A(\encoder1.value[2] ),
    .B(_325_),
    .Y(_326_));
 sky130_fd_sc_hd__nand2_1 _724_ (.A(_324_),
    .B(_326_),
    .Y(_327_));
 sky130_fd_sc_hd__xnor2_1 _725_ (.A(_323_),
    .B(_327_),
    .Y(_328_));
 sky130_fd_sc_hd__nand2_1 _726_ (.A(_315_),
    .B(_328_),
    .Y(_329_));
 sky130_fd_sc_hd__o211a_1 _727_ (.A1(\encoder1.value[2] ),
    .A2(_315_),
    .B1(_329_),
    .C1(_275_),
    .X(_075_));
 sky130_fd_sc_hd__xnor2_1 _728_ (.A(\encoder1.value[3] ),
    .B(_325_),
    .Y(_330_));
 sky130_fd_sc_hd__o21ai_1 _729_ (.A1(_323_),
    .A2(_327_),
    .B1(_326_),
    .Y(_331_));
 sky130_fd_sc_hd__a21bo_1 _730_ (.A1(_330_),
    .A2(_331_),
    .B1_N(_314_),
    .X(_332_));
 sky130_fd_sc_hd__o21bai_1 _731_ (.A1(_330_),
    .A2(_331_),
    .B1_N(_332_),
    .Y(_333_));
 sky130_fd_sc_hd__o211a_1 _732_ (.A1(\encoder1.value[3] ),
    .A2(_315_),
    .B1(_333_),
    .C1(_275_),
    .X(_076_));
 sky130_fd_sc_hd__o21ai_1 _733_ (.A1(\encoder1.value[3] ),
    .A2(\encoder1.value[2] ),
    .B1(_325_),
    .Y(_334_));
 sky130_fd_sc_hd__o31a_1 _734_ (.A1(_323_),
    .A2(_327_),
    .A3(_330_),
    .B1(_334_),
    .X(_335_));
 sky130_fd_sc_hd__xnor2_1 _735_ (.A(\encoder1.value[4] ),
    .B(_325_),
    .Y(_336_));
 sky130_fd_sc_hd__and2_1 _736_ (.A(_335_),
    .B(_336_),
    .X(_337_));
 sky130_fd_sc_hd__nor2_1 _737_ (.A(_335_),
    .B(_336_),
    .Y(_338_));
 sky130_fd_sc_hd__o21ai_1 _738_ (.A1(_337_),
    .A2(_338_),
    .B1(_314_),
    .Y(_339_));
 sky130_fd_sc_hd__o211a_1 _739_ (.A1(\encoder1.value[4] ),
    .A2(_315_),
    .B1(_339_),
    .C1(_275_),
    .X(_077_));
 sky130_fd_sc_hd__xnor2_1 _740_ (.A(\encoder1.value[5] ),
    .B(_325_),
    .Y(_340_));
 sky130_fd_sc_hd__a21o_1 _741_ (.A1(\encoder1.value[4] ),
    .A2(_325_),
    .B1(_338_),
    .X(_341_));
 sky130_fd_sc_hd__nor2_1 _742_ (.A(_340_),
    .B(_341_),
    .Y(_342_));
 sky130_fd_sc_hd__a21bo_1 _743_ (.A1(_340_),
    .A2(_341_),
    .B1_N(_314_),
    .X(_343_));
 sky130_fd_sc_hd__o221a_1 _744_ (.A1(\encoder1.value[5] ),
    .A2(_315_),
    .B1(_342_),
    .B2(_343_),
    .C1(_220_),
    .X(_078_));
 sky130_fd_sc_hd__nor2_1 _745_ (.A(\encoder1.value[6] ),
    .B(_325_),
    .Y(_344_));
 sky130_fd_sc_hd__nand2_1 _746_ (.A(\encoder1.value[6] ),
    .B(_325_),
    .Y(_345_));
 sky130_fd_sc_hd__or2b_1 _747_ (.A(_344_),
    .B_N(_345_),
    .X(_346_));
 sky130_fd_sc_hd__o21ai_1 _748_ (.A1(\encoder1.value[5] ),
    .A2(\encoder1.value[4] ),
    .B1(_325_),
    .Y(_347_));
 sky130_fd_sc_hd__o31a_1 _749_ (.A1(_335_),
    .A2(_336_),
    .A3(_340_),
    .B1(_347_),
    .X(_348_));
 sky130_fd_sc_hd__xnor2_1 _750_ (.A(_346_),
    .B(_348_),
    .Y(_349_));
 sky130_fd_sc_hd__nand2_1 _751_ (.A(_315_),
    .B(_349_),
    .Y(_350_));
 sky130_fd_sc_hd__o211a_1 _752_ (.A1(\encoder1.value[6] ),
    .A2(_315_),
    .B1(_350_),
    .C1(_275_),
    .X(_079_));
 sky130_fd_sc_hd__o21a_1 _753_ (.A1(_344_),
    .A2(_348_),
    .B1(_345_),
    .X(_351_));
 sky130_fd_sc_hd__xnor2_1 _754_ (.A(_129_),
    .B(_325_),
    .Y(_352_));
 sky130_fd_sc_hd__and2_1 _755_ (.A(_351_),
    .B(_352_),
    .X(_353_));
 sky130_fd_sc_hd__o21ai_1 _756_ (.A1(_351_),
    .A2(_352_),
    .B1(_314_),
    .Y(_354_));
 sky130_fd_sc_hd__o221a_1 _757_ (.A1(\encoder1.value[7] ),
    .A2(_315_),
    .B1(_353_),
    .B2(_354_),
    .C1(_220_),
    .X(_080_));
 sky130_fd_sc_hd__and2_1 _758_ (.A(\debounce1_b.debounced ),
    .B(_190_),
    .X(_355_));
 sky130_fd_sc_hd__clkbuf_1 _759_ (.A(_355_),
    .X(_082_));
 sky130_fd_sc_hd__and2b_1 _760_ (.A_N(\debounce2_a.debounced ),
    .B(\debounce2_b.debounced ),
    .X(_356_));
 sky130_fd_sc_hd__and2b_1 _761_ (.A_N(\debounce2_b.debounced ),
    .B(\debounce2_a.debounced ),
    .X(_357_));
 sky130_fd_sc_hd__and2_1 _762_ (.A(\encoder2.old_b ),
    .B(\encoder2.old_a ),
    .X(_358_));
 sky130_fd_sc_hd__nor2_1 _763_ (.A(\encoder2.old_b ),
    .B(\encoder2.old_a ),
    .Y(_359_));
 sky130_fd_sc_hd__o22a_2 _764_ (.A1(_356_),
    .A2(_357_),
    .B1(_358_),
    .B2(_359_),
    .X(_360_));
 sky130_fd_sc_hd__buf_2 _765_ (.A(_360_),
    .X(_361_));
 sky130_fd_sc_hd__a21oi_1 _766_ (.A1(\encoder2.value[0] ),
    .A2(_360_),
    .B1(_242_),
    .Y(_362_));
 sky130_fd_sc_hd__o21a_1 _767_ (.A1(\encoder2.value[0] ),
    .A2(_361_),
    .B1(_362_),
    .X(_083_));
 sky130_fd_sc_hd__o22a_1 _768_ (.A1(_356_),
    .A2(_358_),
    .B1(_359_),
    .B2(_357_),
    .X(_363_));
 sky130_fd_sc_hd__or2_1 _769_ (.A(\encoder2.value[1] ),
    .B(_363_),
    .X(_364_));
 sky130_fd_sc_hd__nand2_1 _770_ (.A(\encoder2.value[1] ),
    .B(_363_),
    .Y(_365_));
 sky130_fd_sc_hd__a21oi_1 _771_ (.A1(_364_),
    .A2(_365_),
    .B1(\encoder2.value[0] ),
    .Y(_366_));
 sky130_fd_sc_hd__and3_1 _772_ (.A(\encoder2.value[0] ),
    .B(_364_),
    .C(_365_),
    .X(_367_));
 sky130_fd_sc_hd__o21ai_1 _773_ (.A1(_366_),
    .A2(_367_),
    .B1(_360_),
    .Y(_368_));
 sky130_fd_sc_hd__o211a_1 _774_ (.A1(\encoder2.value[1] ),
    .A2(_361_),
    .B1(_368_),
    .C1(_220_),
    .X(_084_));
 sky130_fd_sc_hd__a21boi_1 _775_ (.A1(\encoder2.value[0] ),
    .A2(_364_),
    .B1_N(_365_),
    .Y(_369_));
 sky130_fd_sc_hd__or2_1 _776_ (.A(\encoder2.value[2] ),
    .B(_363_),
    .X(_370_));
 sky130_fd_sc_hd__clkbuf_4 _777_ (.A(_363_),
    .X(_371_));
 sky130_fd_sc_hd__nand2_1 _778_ (.A(\encoder2.value[2] ),
    .B(_371_),
    .Y(_372_));
 sky130_fd_sc_hd__nand2_1 _779_ (.A(_370_),
    .B(_372_),
    .Y(_373_));
 sky130_fd_sc_hd__xnor2_1 _780_ (.A(_369_),
    .B(_373_),
    .Y(_374_));
 sky130_fd_sc_hd__nand2_1 _781_ (.A(_361_),
    .B(_374_),
    .Y(_375_));
 sky130_fd_sc_hd__o211a_1 _782_ (.A1(\encoder2.value[2] ),
    .A2(_361_),
    .B1(_375_),
    .C1(_220_),
    .X(_085_));
 sky130_fd_sc_hd__xnor2_1 _783_ (.A(\encoder2.value[3] ),
    .B(_371_),
    .Y(_376_));
 sky130_fd_sc_hd__o21ai_1 _784_ (.A1(_369_),
    .A2(_373_),
    .B1(_372_),
    .Y(_377_));
 sky130_fd_sc_hd__a21bo_1 _785_ (.A1(_376_),
    .A2(_377_),
    .B1_N(_360_),
    .X(_378_));
 sky130_fd_sc_hd__o21bai_1 _786_ (.A1(_376_),
    .A2(_377_),
    .B1_N(_378_),
    .Y(_379_));
 sky130_fd_sc_hd__o211a_1 _787_ (.A1(\encoder2.value[3] ),
    .A2(_361_),
    .B1(_379_),
    .C1(_220_),
    .X(_086_));
 sky130_fd_sc_hd__o21ai_1 _788_ (.A1(\encoder2.value[3] ),
    .A2(\encoder2.value[2] ),
    .B1(_371_),
    .Y(_380_));
 sky130_fd_sc_hd__o31a_1 _789_ (.A1(_369_),
    .A2(_373_),
    .A3(_376_),
    .B1(_380_),
    .X(_381_));
 sky130_fd_sc_hd__xnor2_1 _790_ (.A(\encoder2.value[4] ),
    .B(_371_),
    .Y(_382_));
 sky130_fd_sc_hd__and2_1 _791_ (.A(_381_),
    .B(_382_),
    .X(_383_));
 sky130_fd_sc_hd__nor2_1 _792_ (.A(_381_),
    .B(_382_),
    .Y(_384_));
 sky130_fd_sc_hd__o21ai_1 _793_ (.A1(_383_),
    .A2(_384_),
    .B1(_360_),
    .Y(_385_));
 sky130_fd_sc_hd__o211a_1 _794_ (.A1(\encoder2.value[4] ),
    .A2(_361_),
    .B1(_385_),
    .C1(_220_),
    .X(_087_));
 sky130_fd_sc_hd__xnor2_1 _795_ (.A(\encoder2.value[5] ),
    .B(_371_),
    .Y(_386_));
 sky130_fd_sc_hd__a21oi_1 _796_ (.A1(\encoder2.value[4] ),
    .A2(_371_),
    .B1(_384_),
    .Y(_387_));
 sky130_fd_sc_hd__xnor2_1 _797_ (.A(_386_),
    .B(_387_),
    .Y(_388_));
 sky130_fd_sc_hd__nor2_1 _798_ (.A(\encoder2.value[5] ),
    .B(_360_),
    .Y(_389_));
 sky130_fd_sc_hd__a211oi_1 _799_ (.A1(_361_),
    .A2(_388_),
    .B1(_389_),
    .C1(_145_),
    .Y(_088_));
 sky130_fd_sc_hd__nor2_1 _800_ (.A(\encoder2.value[6] ),
    .B(_371_),
    .Y(_390_));
 sky130_fd_sc_hd__nand2_1 _801_ (.A(\encoder2.value[6] ),
    .B(_371_),
    .Y(_391_));
 sky130_fd_sc_hd__or2b_1 _802_ (.A(_390_),
    .B_N(_391_),
    .X(_392_));
 sky130_fd_sc_hd__o21ai_1 _803_ (.A1(\encoder2.value[5] ),
    .A2(\encoder2.value[4] ),
    .B1(_371_),
    .Y(_393_));
 sky130_fd_sc_hd__o31a_1 _804_ (.A1(_381_),
    .A2(_382_),
    .A3(_386_),
    .B1(_393_),
    .X(_394_));
 sky130_fd_sc_hd__xnor2_1 _805_ (.A(_392_),
    .B(_394_),
    .Y(_395_));
 sky130_fd_sc_hd__nand2_1 _806_ (.A(_361_),
    .B(_395_),
    .Y(_396_));
 sky130_fd_sc_hd__o211a_1 _807_ (.A1(\encoder2.value[6] ),
    .A2(_361_),
    .B1(_396_),
    .C1(_220_),
    .X(_089_));
 sky130_fd_sc_hd__o21a_1 _808_ (.A1(_390_),
    .A2(_394_),
    .B1(_391_),
    .X(_397_));
 sky130_fd_sc_hd__xnor2_1 _809_ (.A(_146_),
    .B(_371_),
    .Y(_398_));
 sky130_fd_sc_hd__and2_1 _810_ (.A(_397_),
    .B(_398_),
    .X(_399_));
 sky130_fd_sc_hd__o21ai_1 _811_ (.A1(_397_),
    .A2(_398_),
    .B1(_360_),
    .Y(_400_));
 sky130_fd_sc_hd__o221a_1 _812_ (.A1(\encoder2.value[7] ),
    .A2(_361_),
    .B1(_399_),
    .B2(_400_),
    .C1(_220_),
    .X(_090_));
 sky130_fd_sc_hd__and2_1 _813_ (.A(\debounce2_b.debounced ),
    .B(_232_),
    .X(_401_));
 sky130_fd_sc_hd__clkbuf_1 _814_ (.A(_401_),
    .X(_091_));
 sky130_fd_sc_hd__nor2_1 _815_ (.A(_145_),
    .B(\pwm0.count[0] ),
    .Y(_092_));
 sky130_fd_sc_hd__a21o_1 _816_ (.A1(\pwm0.count[1] ),
    .A2(\pwm0.count[0] ),
    .B1(net7),
    .X(_402_));
 sky130_fd_sc_hd__a21oi_1 _817_ (.A1(_117_),
    .A2(_119_),
    .B1(_402_),
    .Y(_093_));
 sky130_fd_sc_hd__a21oi_1 _818_ (.A1(\pwm0.count[1] ),
    .A2(\pwm0.count[0] ),
    .B1(\pwm0.count[2] ),
    .Y(_403_));
 sky130_fd_sc_hd__and3_1 _819_ (.A(\pwm0.count[2] ),
    .B(\pwm0.count[1] ),
    .C(\pwm0.count[0] ),
    .X(_404_));
 sky130_fd_sc_hd__nor3_1 _820_ (.A(_145_),
    .B(_403_),
    .C(_404_),
    .Y(_094_));
 sky130_fd_sc_hd__and2_1 _821_ (.A(\pwm0.count[3] ),
    .B(_404_),
    .X(_405_));
 sky130_fd_sc_hd__o21ai_1 _822_ (.A1(\pwm0.count[3] ),
    .A2(_404_),
    .B1(_162_),
    .Y(_406_));
 sky130_fd_sc_hd__nor2_1 _823_ (.A(_405_),
    .B(_406_),
    .Y(_095_));
 sky130_fd_sc_hd__and3_1 _824_ (.A(\pwm0.count[4] ),
    .B(\pwm0.count[3] ),
    .C(_404_),
    .X(_407_));
 sky130_fd_sc_hd__o21ai_1 _825_ (.A1(\pwm0.count[4] ),
    .A2(_405_),
    .B1(_162_),
    .Y(_408_));
 sky130_fd_sc_hd__nor2_1 _826_ (.A(_407_),
    .B(_408_),
    .Y(_096_));
 sky130_fd_sc_hd__and2_1 _827_ (.A(\pwm0.count[5] ),
    .B(_407_),
    .X(_409_));
 sky130_fd_sc_hd__nor2_1 _828_ (.A(_242_),
    .B(_409_),
    .Y(_410_));
 sky130_fd_sc_hd__o21a_1 _829_ (.A1(\pwm0.count[5] ),
    .A2(_407_),
    .B1(_410_),
    .X(_097_));
 sky130_fd_sc_hd__and3_1 _830_ (.A(\pwm0.count[6] ),
    .B(\pwm0.count[5] ),
    .C(_407_),
    .X(_411_));
 sky130_fd_sc_hd__o21ai_1 _831_ (.A1(\pwm0.count[6] ),
    .A2(_409_),
    .B1(_162_),
    .Y(_412_));
 sky130_fd_sc_hd__nor2_1 _832_ (.A(_411_),
    .B(_412_),
    .Y(_098_));
 sky130_fd_sc_hd__a21oi_1 _833_ (.A1(\pwm0.count[7] ),
    .A2(_411_),
    .B1(_242_),
    .Y(_413_));
 sky130_fd_sc_hd__o21a_1 _834_ (.A1(\pwm0.count[7] ),
    .A2(_411_),
    .B1(_413_),
    .X(_099_));
 sky130_fd_sc_hd__nor2_1 _835_ (.A(_145_),
    .B(\pwm1.count[0] ),
    .Y(_100_));
 sky130_fd_sc_hd__a21oi_1 _836_ (.A1(\pwm1.count[1] ),
    .A2(\pwm1.count[0] ),
    .B1(_242_),
    .Y(_414_));
 sky130_fd_sc_hd__o21a_1 _837_ (.A1(\pwm1.count[1] ),
    .A2(\pwm1.count[0] ),
    .B1(_414_),
    .X(_101_));
 sky130_fd_sc_hd__a21oi_1 _838_ (.A1(\pwm1.count[1] ),
    .A2(\pwm1.count[0] ),
    .B1(\pwm1.count[2] ),
    .Y(_415_));
 sky130_fd_sc_hd__and3_1 _839_ (.A(\pwm1.count[2] ),
    .B(\pwm1.count[1] ),
    .C(\pwm1.count[0] ),
    .X(_416_));
 sky130_fd_sc_hd__nor3_1 _840_ (.A(_145_),
    .B(_415_),
    .C(_416_),
    .Y(_102_));
 sky130_fd_sc_hd__and2_1 _841_ (.A(\pwm1.count[3] ),
    .B(_416_),
    .X(_417_));
 sky130_fd_sc_hd__o21ai_1 _842_ (.A1(\pwm1.count[3] ),
    .A2(_416_),
    .B1(_162_),
    .Y(_418_));
 sky130_fd_sc_hd__nor2_1 _843_ (.A(_417_),
    .B(_418_),
    .Y(_103_));
 sky130_fd_sc_hd__and3_1 _844_ (.A(\pwm1.count[4] ),
    .B(\pwm1.count[3] ),
    .C(_416_),
    .X(_419_));
 sky130_fd_sc_hd__o21ai_1 _845_ (.A1(\pwm1.count[4] ),
    .A2(_417_),
    .B1(_169_),
    .Y(_420_));
 sky130_fd_sc_hd__nor2_1 _846_ (.A(_419_),
    .B(_420_),
    .Y(_104_));
 sky130_fd_sc_hd__and2_1 _847_ (.A(\pwm1.count[5] ),
    .B(_419_),
    .X(_421_));
 sky130_fd_sc_hd__nor2_1 _848_ (.A(net7),
    .B(_421_),
    .Y(_422_));
 sky130_fd_sc_hd__o21a_1 _849_ (.A1(\pwm1.count[5] ),
    .A2(_419_),
    .B1(_422_),
    .X(_105_));
 sky130_fd_sc_hd__and3_1 _850_ (.A(\pwm1.count[6] ),
    .B(\pwm1.count[5] ),
    .C(_419_),
    .X(_423_));
 sky130_fd_sc_hd__o21ai_1 _851_ (.A1(\pwm1.count[6] ),
    .A2(_421_),
    .B1(_169_),
    .Y(_424_));
 sky130_fd_sc_hd__nor2_1 _852_ (.A(_423_),
    .B(_424_),
    .Y(_106_));
 sky130_fd_sc_hd__a21oi_1 _853_ (.A1(\pwm1.count[7] ),
    .A2(_423_),
    .B1(_242_),
    .Y(_425_));
 sky130_fd_sc_hd__o21a_1 _854_ (.A1(\pwm1.count[7] ),
    .A2(_423_),
    .B1(_425_),
    .X(_107_));
 sky130_fd_sc_hd__dfxtp_1 _855_ (.CLK(clknet_3_6__leaf_clk),
    .D(_000_),
    .Q(\debounce0_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _856_ (.CLK(clknet_3_6__leaf_clk),
    .D(_001_),
    .Q(\debounce0_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _857_ (.CLK(clknet_3_6__leaf_clk),
    .D(_002_),
    .Q(\debounce0_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _858_ (.CLK(clknet_3_6__leaf_clk),
    .D(_003_),
    .Q(\debounce0_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _859_ (.CLK(clknet_3_7__leaf_clk),
    .D(_004_),
    .Q(\debounce0_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _860_ (.CLK(clknet_3_7__leaf_clk),
    .D(_005_),
    .Q(\debounce0_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _861_ (.CLK(clknet_3_7__leaf_clk),
    .D(_006_),
    .Q(\debounce0_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _862_ (.CLK(clknet_3_7__leaf_clk),
    .D(_007_),
    .Q(\debounce0_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _863_ (.CLK(clknet_3_7__leaf_clk),
    .D(_008_),
    .Q(\debounce0_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _864_ (.CLK(clknet_3_7__leaf_clk),
    .D(_009_),
    .Q(\debounce0_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _865_ (.CLK(clknet_3_7__leaf_clk),
    .D(_010_),
    .Q(\debounce0_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _866_ (.CLK(clknet_3_7__leaf_clk),
    .D(_011_),
    .Q(\debounce0_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _867_ (.CLK(clknet_3_7__leaf_clk),
    .D(_012_),
    .Q(\debounce0_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _868_ (.CLK(clknet_3_7__leaf_clk),
    .D(_013_),
    .Q(\debounce0_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _869_ (.CLK(clknet_3_7__leaf_clk),
    .D(_014_),
    .Q(\debounce0_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _870_ (.CLK(clknet_3_7__leaf_clk),
    .D(_015_),
    .Q(\debounce0_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _871_ (.CLK(clknet_3_7__leaf_clk),
    .D(_016_),
    .Q(\debounce0_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _872_ (.CLK(clknet_3_7__leaf_clk),
    .D(_017_),
    .Q(\debounce0_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _873_ (.CLK(clknet_3_5__leaf_clk),
    .D(_018_),
    .Q(\debounce1_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _874_ (.CLK(clknet_3_5__leaf_clk),
    .D(_019_),
    .Q(\debounce1_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _875_ (.CLK(clknet_3_5__leaf_clk),
    .D(_020_),
    .Q(\debounce1_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _876_ (.CLK(clknet_3_5__leaf_clk),
    .D(_021_),
    .Q(\debounce1_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _877_ (.CLK(clknet_3_5__leaf_clk),
    .D(_022_),
    .Q(\debounce1_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _878_ (.CLK(clknet_3_5__leaf_clk),
    .D(_023_),
    .Q(\debounce1_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _879_ (.CLK(clknet_3_5__leaf_clk),
    .D(_024_),
    .Q(\debounce1_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _880_ (.CLK(clknet_3_5__leaf_clk),
    .D(_025_),
    .Q(\debounce1_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _881_ (.CLK(clknet_3_5__leaf_clk),
    .D(_026_),
    .Q(\debounce1_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _882_ (.CLK(clknet_3_6__leaf_clk),
    .D(_027_),
    .Q(\debounce1_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _883_ (.CLK(clknet_3_6__leaf_clk),
    .D(_028_),
    .Q(\debounce1_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _884_ (.CLK(clknet_3_7__leaf_clk),
    .D(_029_),
    .Q(\debounce1_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _885_ (.CLK(clknet_3_6__leaf_clk),
    .D(_030_),
    .Q(\debounce1_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _886_ (.CLK(clknet_3_6__leaf_clk),
    .D(_031_),
    .Q(\debounce1_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _887_ (.CLK(clknet_3_7__leaf_clk),
    .D(_032_),
    .Q(\debounce1_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _888_ (.CLK(clknet_3_7__leaf_clk),
    .D(_033_),
    .Q(\debounce1_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _889_ (.CLK(clknet_3_5__leaf_clk),
    .D(_034_),
    .Q(\debounce1_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _890_ (.CLK(clknet_3_5__leaf_clk),
    .D(_035_),
    .Q(\debounce1_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _891_ (.CLK(clknet_3_1__leaf_clk),
    .D(_036_),
    .Q(\debounce2_a.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _892_ (.CLK(clknet_3_1__leaf_clk),
    .D(_037_),
    .Q(\debounce2_a.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _893_ (.CLK(clknet_3_1__leaf_clk),
    .D(_038_),
    .Q(\debounce2_a.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _894_ (.CLK(clknet_3_1__leaf_clk),
    .D(_039_),
    .Q(\debounce2_a.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _895_ (.CLK(clknet_3_1__leaf_clk),
    .D(_040_),
    .Q(\debounce2_a.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _896_ (.CLK(clknet_3_4__leaf_clk),
    .D(_041_),
    .Q(\debounce2_a.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _897_ (.CLK(clknet_3_4__leaf_clk),
    .D(_042_),
    .Q(\debounce2_a.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _898_ (.CLK(clknet_3_1__leaf_clk),
    .D(_043_),
    .Q(\debounce2_a.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _899_ (.CLK(clknet_3_1__leaf_clk),
    .D(_044_),
    .Q(\debounce2_a.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _900_ (.CLK(clknet_3_4__leaf_clk),
    .D(_045_),
    .Q(\debounce2_b.debounced ));
 sky130_fd_sc_hd__dfxtp_1 _901_ (.CLK(clknet_3_0__leaf_clk),
    .D(_046_),
    .Q(\pwm2.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _902_ (.CLK(clknet_3_0__leaf_clk),
    .D(_047_),
    .Q(\pwm2.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _903_ (.CLK(clknet_3_2__leaf_clk),
    .D(_048_),
    .Q(\pwm2.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _904_ (.CLK(clknet_3_3__leaf_clk),
    .D(_049_),
    .Q(\pwm2.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _905_ (.CLK(clknet_3_2__leaf_clk),
    .D(_050_),
    .Q(\pwm2.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _906_ (.CLK(clknet_3_2__leaf_clk),
    .D(_051_),
    .Q(\pwm2.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _907_ (.CLK(clknet_3_2__leaf_clk),
    .D(_052_),
    .Q(\pwm2.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _908_ (.CLK(clknet_3_2__leaf_clk),
    .D(_053_),
    .Q(\pwm2.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _909_ (.CLK(clknet_3_7__leaf_clk),
    .D(_054_),
    .Q(\encoder0.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _910_ (.CLK(clknet_3_4__leaf_clk),
    .D(_055_),
    .Q(\debounce2_b.button_hist[0] ));
 sky130_fd_sc_hd__dfxtp_1 _911_ (.CLK(clknet_3_5__leaf_clk),
    .D(_056_),
    .Q(\debounce2_b.button_hist[1] ));
 sky130_fd_sc_hd__dfxtp_1 _912_ (.CLK(clknet_3_5__leaf_clk),
    .D(_057_),
    .Q(\debounce2_b.button_hist[2] ));
 sky130_fd_sc_hd__dfxtp_1 _913_ (.CLK(clknet_3_4__leaf_clk),
    .D(_058_),
    .Q(\debounce2_b.button_hist[3] ));
 sky130_fd_sc_hd__dfxtp_1 _914_ (.CLK(clknet_3_4__leaf_clk),
    .D(_059_),
    .Q(\debounce2_b.button_hist[4] ));
 sky130_fd_sc_hd__dfxtp_1 _915_ (.CLK(clknet_3_4__leaf_clk),
    .D(_060_),
    .Q(\debounce2_b.button_hist[5] ));
 sky130_fd_sc_hd__dfxtp_1 _916_ (.CLK(clknet_3_4__leaf_clk),
    .D(_061_),
    .Q(\debounce2_b.button_hist[6] ));
 sky130_fd_sc_hd__dfxtp_1 _917_ (.CLK(clknet_3_5__leaf_clk),
    .D(_062_),
    .Q(\debounce2_b.button_hist[7] ));
 sky130_fd_sc_hd__dfxtp_1 _918_ (.CLK(clknet_3_6__leaf_clk),
    .D(_063_),
    .Q(\encoder0.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _919_ (.CLK(clknet_3_6__leaf_clk),
    .D(_064_),
    .Q(\encoder0.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _920_ (.CLK(clknet_3_3__leaf_clk),
    .D(_065_),
    .Q(\encoder0.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _921_ (.CLK(clknet_3_3__leaf_clk),
    .D(_066_),
    .Q(\encoder0.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _922_ (.CLK(clknet_3_2__leaf_clk),
    .D(_067_),
    .Q(\encoder0.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _923_ (.CLK(clknet_3_2__leaf_clk),
    .D(_068_),
    .Q(\encoder0.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _924_ (.CLK(clknet_3_3__leaf_clk),
    .D(_069_),
    .Q(\encoder0.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _925_ (.CLK(clknet_3_6__leaf_clk),
    .D(_070_),
    .Q(\encoder0.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _926_ (.CLK(clknet_3_5__leaf_clk),
    .D(_071_),
    .Q(\encoder1.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _927_ (.CLK(clknet_3_6__leaf_clk),
    .D(_072_),
    .Q(\encoder0.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _928_ (.CLK(clknet_3_1__leaf_clk),
    .D(_073_),
    .Q(\encoder1.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _929_ (.CLK(clknet_3_4__leaf_clk),
    .D(_074_),
    .Q(\encoder1.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _930_ (.CLK(clknet_3_4__leaf_clk),
    .D(_075_),
    .Q(\encoder1.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _931_ (.CLK(clknet_3_1__leaf_clk),
    .D(_076_),
    .Q(\encoder1.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _932_ (.CLK(clknet_3_1__leaf_clk),
    .D(_077_),
    .Q(\encoder1.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _933_ (.CLK(clknet_3_0__leaf_clk),
    .D(_078_),
    .Q(\encoder1.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _934_ (.CLK(clknet_3_0__leaf_clk),
    .D(_079_),
    .Q(\encoder1.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _935_ (.CLK(clknet_3_0__leaf_clk),
    .D(_080_),
    .Q(\encoder1.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _936_ (.CLK(clknet_3_6__leaf_clk),
    .D(_081_),
    .Q(\encoder2.old_a ));
 sky130_fd_sc_hd__dfxtp_1 _937_ (.CLK(clknet_3_4__leaf_clk),
    .D(_082_),
    .Q(\encoder1.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _938_ (.CLK(clknet_3_0__leaf_clk),
    .D(_083_),
    .Q(\encoder2.value[0] ));
 sky130_fd_sc_hd__dfxtp_1 _939_ (.CLK(clknet_3_0__leaf_clk),
    .D(_084_),
    .Q(\encoder2.value[1] ));
 sky130_fd_sc_hd__dfxtp_1 _940_ (.CLK(clknet_3_2__leaf_clk),
    .D(_085_),
    .Q(\encoder2.value[2] ));
 sky130_fd_sc_hd__dfxtp_1 _941_ (.CLK(clknet_3_2__leaf_clk),
    .D(_086_),
    .Q(\encoder2.value[3] ));
 sky130_fd_sc_hd__dfxtp_1 _942_ (.CLK(clknet_3_2__leaf_clk),
    .D(_087_),
    .Q(\encoder2.value[4] ));
 sky130_fd_sc_hd__dfxtp_1 _943_ (.CLK(clknet_3_2__leaf_clk),
    .D(_088_),
    .Q(\encoder2.value[5] ));
 sky130_fd_sc_hd__dfxtp_1 _944_ (.CLK(clknet_3_2__leaf_clk),
    .D(_089_),
    .Q(\encoder2.value[6] ));
 sky130_fd_sc_hd__dfxtp_1 _945_ (.CLK(clknet_3_2__leaf_clk),
    .D(_090_),
    .Q(\encoder2.value[7] ));
 sky130_fd_sc_hd__dfxtp_1 _946_ (.CLK(clknet_3_0__leaf_clk),
    .D(_091_),
    .Q(\encoder2.old_b ));
 sky130_fd_sc_hd__dfxtp_1 _947_ (.CLK(clknet_3_3__leaf_clk),
    .D(_092_),
    .Q(\pwm0.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _948_ (.CLK(clknet_3_3__leaf_clk),
    .D(_093_),
    .Q(\pwm0.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _949_ (.CLK(clknet_3_3__leaf_clk),
    .D(_094_),
    .Q(\pwm0.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _950_ (.CLK(clknet_3_3__leaf_clk),
    .D(_095_),
    .Q(\pwm0.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _951_ (.CLK(clknet_3_3__leaf_clk),
    .D(_096_),
    .Q(\pwm0.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _952_ (.CLK(clknet_3_6__leaf_clk),
    .D(_097_),
    .Q(\pwm0.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _953_ (.CLK(clknet_3_6__leaf_clk),
    .D(_098_),
    .Q(\pwm0.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _954_ (.CLK(clknet_3_6__leaf_clk),
    .D(_099_),
    .Q(\pwm0.count[7] ));
 sky130_fd_sc_hd__dfxtp_1 _955_ (.CLK(clknet_3_0__leaf_clk),
    .D(_100_),
    .Q(\pwm1.count[0] ));
 sky130_fd_sc_hd__dfxtp_1 _956_ (.CLK(clknet_3_1__leaf_clk),
    .D(_101_),
    .Q(\pwm1.count[1] ));
 sky130_fd_sc_hd__dfxtp_1 _957_ (.CLK(clknet_3_0__leaf_clk),
    .D(_102_),
    .Q(\pwm1.count[2] ));
 sky130_fd_sc_hd__dfxtp_1 _958_ (.CLK(clknet_3_0__leaf_clk),
    .D(_103_),
    .Q(\pwm1.count[3] ));
 sky130_fd_sc_hd__dfxtp_1 _959_ (.CLK(clknet_3_0__leaf_clk),
    .D(_104_),
    .Q(\pwm1.count[4] ));
 sky130_fd_sc_hd__dfxtp_1 _960_ (.CLK(clknet_3_0__leaf_clk),
    .D(_105_),
    .Q(\pwm1.count[5] ));
 sky130_fd_sc_hd__dfxtp_1 _961_ (.CLK(clknet_3_0__leaf_clk),
    .D(_106_),
    .Q(\pwm1.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 _962_ (.CLK(clknet_3_0__leaf_clk),
    .D(_107_),
    .Q(\pwm1.count[7] ));
 sky130_fd_sc_hd__conb_1 rgb_mixer_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 rgb_mixer_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 rgb_mixer_15 (.LO(net15));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_1 _967_ (.A(net7),
    .X(net11));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(enc0_a),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(enc0_b),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(enc1_a),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(enc1_b),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(enc2_a),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(enc2_b),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_4 input7 (.A(reset),
    .X(net7));
 sky130_fd_sc_hd__buf_2 output8 (.A(net8),
    .X(pwm0_out));
 sky130_fd_sc_hd__buf_2 output9 (.A(net9),
    .X(pwm1_out));
 sky130_fd_sc_hd__buf_2 output10 (.A(net10),
    .X(pwm2_out));
 sky130_fd_sc_hd__buf_2 output11 (.A(net11),
    .X(sync));
 sky130_fd_sc_hd__conb_1 rgb_mixer_12 (.LO(net12));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(net5));
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_32 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_227 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_219 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_232 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_294 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_392 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_287 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_234 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_352 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_224 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_405 ();
 assign io_oeb[0] = net12;
 assign io_oeb[1] = net13;
 assign io_oeb[2] = net14;
 assign io_oeb[3] = net15;
endmodule

